--------------------------------------------------------------------------------
-- saa5050_rom_data.vhd                                                       --
-- Character ROM for the SAA5050.                                             --
--------------------------------------------------------------------------------
-- (C) Copyright 2022 Adam Barnes <ambarnes@gmail.com>                        --
-- This file is part of The Tyto Project. The Tyto Project is free software:  --
-- you can redistribute it and/or modify it under the terms of the GNU Lesser --
-- General Public License as published by the Free Software Foundation,       --
-- either version 3 of the License, or (at your option) any later version.    --
-- The Tyto Project is distributed in the hope that it will be useful, but    --
-- WITHOUT ANY WARRANTY; without even the implied warranty of MERCHANTABILITY --
-- or FITNESS FOR A PARTICULAR PURPOSE. See the GNU Lesser General Public     --
-- License for more details. You should have received a copy of the GNU       --
-- Lesser General Public License along with The Tyto Project. If not, see     --
-- https://www.gnu.org/licenses/.                                             --
--------------------------------------------------------------------------------

-- Original teletext character set = 96 characters, each 9 (v) x 5 (h) pixels.
-- These are padded with empty pixels to 6 by 10, and a clever rounding feature
-- doubles the displayed resolution to 12 x 20.
-- Each character is stored in ROM as 16 words (v) x 5 bits (h)
-- 96 characters + 32 spare = 128; 128 x 16 x 8 bits = 16kBits/2kbytes total

library ieee;
use ieee.std_logic_1164.all;

package saa5050_rom_data_pkg is

    type rom_data_t is array(0 to 2047) of std_logic_vector(4 downto 0);
    constant rom_data : rom_data_t := (
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00100",
        "00100",
        "00100",
        "00100",
        "00100",
        "00000",
        "00100",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "01010",
        "01010",
        "01010",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00110",
        "01000",
        "01000",
        "11100",
        "01000",
        "01000",
        "11111",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "01110",
        "10101",
        "10100",
        "01110",
        "00101",
        "10101",
        "01110",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "11000",
        "11001",
        "00010",
        "00100",
        "01000",
        "10011",
        "00011",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "01000",
        "10100",
        "10100",
        "01000",
        "10101",
        "10010",
        "01101",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00100",
        "00100",
        "00100",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00010",
        "00100",
        "01000",
        "01000",
        "01000",
        "00100",
        "00010",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "01000",
        "00100",
        "00010",
        "00010",
        "00010",
        "00100",
        "01000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00100",
        "10101",
        "01110",
        "00100",
        "01110",
        "10101",
        "00100",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00100",
        "00100",
        "11111",
        "00100",
        "00100",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00100",
        "00100",
        "01000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "01110",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00100",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00001",
        "00010",
        "00100",
        "01000",
        "10000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00100",
        "01010",
        "10001",
        "10001",
        "10001",
        "01010",
        "00100",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00100",
        "01100",
        "00100",
        "00100",
        "00100",
        "00100",
        "01110",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "01110",
        "10001",
        "00001",
        "00110",
        "01000",
        "10000",
        "11111",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "11111",
        "00001",
        "00010",
        "00110",
        "00001",
        "10001",
        "01110",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00010",
        "00110",
        "01010",
        "10010",
        "11111",
        "00010",
        "00010",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "11111",
        "10000",
        "11110",
        "00001",
        "00001",
        "10001",
        "01110",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00110",
        "01000",
        "10000",
        "11110",
        "10001",
        "10001",
        "01110",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "11111",
        "00001",
        "00010",
        "00100",
        "01000",
        "01000",
        "01000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "01110",
        "10001",
        "10001",
        "01110",
        "10001",
        "10001",
        "01110",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "01110",
        "10001",
        "10001",
        "01111",
        "00001",
        "00010",
        "01100",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00100",
        "00000",
        "00000",
        "00000",
        "00100",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00100",
        "00000",
        "00000",
        "00100",
        "00100",
        "01000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00010",
        "00100",
        "01000",
        "10000",
        "01000",
        "00100",
        "00010",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "11111",
        "00000",
        "11111",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "01000",
        "00100",
        "00010",
        "00001",
        "00010",
        "00100",
        "01000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "01110",
        "10001",
        "00010",
        "00100",
        "00100",
        "00000",
        "00100",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "01110",
        "10001",
        "10111",
        "10101",
        "10111",
        "10000",
        "01110",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00100",
        "01010",
        "10001",
        "10001",
        "11111",
        "10001",
        "10001",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "11110",
        "10001",
        "10001",
        "11110",
        "10001",
        "10001",
        "11110",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "01110",
        "10001",
        "10000",
        "10000",
        "10000",
        "10001",
        "01110",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "11110",
        "10001",
        "10001",
        "10001",
        "10001",
        "10001",
        "11110",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "11111",
        "10000",
        "10000",
        "11110",
        "10000",
        "10000",
        "11111",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "11111",
        "10000",
        "10000",
        "11110",
        "10000",
        "10000",
        "10000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "01110",
        "10001",
        "10000",
        "10000",
        "10011",
        "10001",
        "01110",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "10001",
        "10001",
        "10001",
        "11111",
        "10001",
        "10001",
        "10001",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "01110",
        "00100",
        "00100",
        "00100",
        "00100",
        "00100",
        "01110",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00001",
        "00001",
        "00001",
        "00001",
        "00001",
        "10001",
        "01110",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "10001",
        "10010",
        "10100",
        "11000",
        "10100",
        "10010",
        "10001",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "10000",
        "10000",
        "10000",
        "10000",
        "10000",
        "10000",
        "11111",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "10001",
        "11011",
        "10101",
        "10101",
        "10001",
        "10001",
        "10001",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "10001",
        "10001",
        "11001",
        "10101",
        "10011",
        "10001",
        "10001",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "01110",
        "10001",
        "10001",
        "10001",
        "10001",
        "10001",
        "01110",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "11110",
        "10001",
        "10001",
        "11110",
        "10000",
        "10000",
        "10000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "01110",
        "10001",
        "10001",
        "10001",
        "10101",
        "10010",
        "01101",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "11110",
        "10001",
        "10001",
        "11110",
        "10100",
        "10010",
        "10001",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "01110",
        "10001",
        "10000",
        "01110",
        "00001",
        "10001",
        "01110",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "11111",
        "00100",
        "00100",
        "00100",
        "00100",
        "00100",
        "00100",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "10001",
        "10001",
        "10001",
        "10001",
        "10001",
        "10001",
        "01110",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "10001",
        "10001",
        "10001",
        "01010",
        "01010",
        "00100",
        "00100",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "10001",
        "10001",
        "10001",
        "10101",
        "10101",
        "10101",
        "01010",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "10001",
        "10001",
        "01010",
        "00100",
        "01010",
        "10001",
        "10001",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "10001",
        "10001",
        "01010",
        "00100",
        "00100",
        "00100",
        "00100",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "11111",
        "00001",
        "00010",
        "00100",
        "01000",
        "10000",
        "11111",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00100",
        "01000",
        "11111",
        "01000",
        "00100",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "10000",
        "10000",
        "10000",
        "10110",
        "00001",
        "00010",
        "00100",
        "00111",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00100",
        "00010",
        "11111",
        "00010",
        "00100",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00100",
        "01110",
        "10101",
        "00100",
        "00100",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "01010",
        "01010",
        "11111",
        "01010",
        "11111",
        "01010",
        "01010",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "11111",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "01110",
        "00001",
        "01111",
        "10001",
        "01111",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "10000",
        "10000",
        "11110",
        "10001",
        "10001",
        "10001",
        "11110",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "01111",
        "10000",
        "10000",
        "10000",
        "01111",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00001",
        "00001",
        "01111",
        "10001",
        "10001",
        "10001",
        "01111",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "01110",
        "10001",
        "11111",
        "10000",
        "01110",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00010",
        "00100",
        "00100",
        "01110",
        "00100",
        "00100",
        "00100",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "01111",
        "10001",
        "10001",
        "10001",
        "01111",
        "00001",
        "01110",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "10000",
        "10000",
        "11110",
        "10001",
        "10001",
        "10001",
        "10001",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00100",
        "00000",
        "01100",
        "00100",
        "00100",
        "00100",
        "01110",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00100",
        "00000",
        "00100",
        "00100",
        "00100",
        "00100",
        "00100",
        "00100",
        "01000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "01000",
        "01000",
        "01001",
        "01010",
        "01100",
        "01010",
        "01001",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "01100",
        "00100",
        "00100",
        "00100",
        "00100",
        "00100",
        "01110",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "11010",
        "10101",
        "10101",
        "10101",
        "10101",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "11110",
        "10001",
        "10001",
        "10001",
        "10001",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "01110",
        "10001",
        "10001",
        "10001",
        "01110",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "11110",
        "10001",
        "10001",
        "10001",
        "11110",
        "10000",
        "10000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "01111",
        "10001",
        "10001",
        "10001",
        "01111",
        "00001",
        "00001",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "01011",
        "01100",
        "01000",
        "01000",
        "01000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "01111",
        "10000",
        "01110",
        "00001",
        "11110",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00100",
        "00100",
        "01110",
        "00100",
        "00100",
        "00100",
        "00010",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "10001",
        "10001",
        "10001",
        "10001",
        "01111",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "10001",
        "10001",
        "01010",
        "01010",
        "00100",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "10001",
        "10001",
        "10101",
        "10101",
        "01010",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "10001",
        "01010",
        "00100",
        "01010",
        "10001",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "10001",
        "10001",
        "10001",
        "10001",
        "01111",
        "00001",
        "01110",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "11111",
        "00010",
        "00100",
        "01000",
        "11111",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "01000",
        "01000",
        "01000",
        "01001",
        "00011",
        "00101",
        "00111",
        "00001",
        "00001",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "01010",
        "01010",
        "01010",
        "01010",
        "01010",
        "01010",
        "01010",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "11000",
        "00100",
        "11000",
        "00100",
        "11001",
        "00011",
        "00101",
        "00111",
        "00001",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00100",
        "00000",
        "11111",
        "00000",
        "00100",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "11111",
        "11111",
        "11111",
        "11111",
        "11111",
        "11111",
        "11111",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000",
        "00000"
    );

end package saa5050_rom_data_pkg;
