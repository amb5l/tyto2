--------------------------------------------------------------------------------
-- tb_hdmi_tpg_mega65_r5.vhd                                                  --
-- Simulation testbench for hdmi_tpg_mega65_r5.vhd.                           --
--------------------------------------------------------------------------------
-- (C) Copyright 2024 Adam Barnes <ambarnes@gmail.com>                        --
-- This file is part of The Tyto Project. The Tyto Project is free software:  --
-- you can redistribute it and/or modify it under the terms of the GNU Lesser --
-- General Public License as published by the Free Software Foundation,       --
-- either version 3 of the License, or (at your option) any later version.    --
-- The Tyto Project is distributed in the hope that it will be useful, but    --
-- WITHOUT ANY WARRANTY; without even the implied warranty of MERCHANTABILITY --
-- or FITNESS FOR A PARTICULAR PURPOSE. See the GNU Lesser General Public     --
-- License for more details. You should have received a copy of the GNU       --
-- Lesser General Public License along with The Tyto Project. If not, see     --
-- https://www.gnu.org/licenses/.                                             --
--------------------------------------------------------------------------------

entity tb_hdmi_tpg_mega65_r5 is
end entity tb_hdmi_tpg_mega65_r5;

architecture sim of tb_hdmi_tpg_mega65_r5 is
begin
end architecture sim;
