entity test_fit_hram_ctrl is
end entity test_fit_hram_ctrl;

architecture rtl of test_fit_hram_ctrl is

begin

  CTRL: component hram_ctrl
    generic map (

    )
    port map (

    );

end architecture rtl;
