package OsvvmTestCommonPkg is
  constant OSVVM_RESULTS_DIR   : string := "" ;
end package OsvvmTestCommonPkg ;
