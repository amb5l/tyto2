package OsvvmTestCommonPkg is
  constant OSVVM_RESULTS_DIR   : string := "" ;
  --constant OSVVM_PATH_TO_TESTS : string := "../../OsvvmLibraries/" ;
end package OsvvmTestCommonPkg ; 
