library ieee;
use ieee.std_logic_1164.all;

package char_rom_437_8x16_pkg is

    component char_rom_437_8x16 is
        port (
            clk : in    std_logic;
            r   : in    std_logic_vector(3 downto 0);
            a   : in    std_logic_vector(7 downto 0);
            d   : out   std_logic_vector(7 downto 0)
        );
    end component char_rom_437_8x16;

end package char_rom_437_8x16_pkg;

library ieee;
use ieee.std_logic_1164.all;

entity char_rom_437_8x16 is
    port (
        clk : in    std_logic;
        r   : in    std_logic_vector(3 downto 0);
        a   : in    std_logic_vector(7 downto 0);
        d   : out   std_logic_vector(7 downto 0)
    );
end entity char_rom_437_8x16;

architecture behavioural of char_rom_437_8x16 is
begin

    process(clk)
    begin
        if rising_edge(clk) then
            case a & r is

                when x"00" & "0000" => d <= "00000000"; -- ........
                when x"00" & "0001" => d <= "00000000"; -- ........
                when x"00" & "0010" => d <= "00000000"; -- ........
                when x"00" & "0011" => d <= "00000000"; -- ........
                when x"00" & "0100" => d <= "00000000"; -- ........
                when x"00" & "0101" => d <= "00000000"; -- ........
                when x"00" & "0110" => d <= "00000000"; -- ........
                when x"00" & "0111" => d <= "00000000"; -- ........
                when x"00" & "1000" => d <= "00000000"; -- ........
                when x"00" & "1001" => d <= "00000000"; -- ........
                when x"00" & "1010" => d <= "00000000"; -- ........
                when x"00" & "1011" => d <= "00000000"; -- ........
                when x"00" & "1100" => d <= "00000000"; -- ........
                when x"00" & "1101" => d <= "00000000"; -- ........
                when x"00" & "1110" => d <= "00000000"; -- ........
                when x"00" & "1111" => d <= "00000000"; -- ........

                when x"01" & "0000" => d <= "00000000"; -- ........
                when x"01" & "0001" => d <= "00000000"; -- ........
                when x"01" & "0010" => d <= "01111110"; -- .######.
                when x"01" & "0011" => d <= "10000001"; -- #......#
                when x"01" & "0100" => d <= "10100101"; -- #.#..#.#
                when x"01" & "0101" => d <= "10000001"; -- #......#
                when x"01" & "0110" => d <= "10000001"; -- #......#
                when x"01" & "0111" => d <= "10111101"; -- #.####.#
                when x"01" & "1000" => d <= "10011001"; -- #..##..#
                when x"01" & "1001" => d <= "10000001"; -- #......#
                when x"01" & "1010" => d <= "10000001"; -- #......#
                when x"01" & "1011" => d <= "01111110"; -- .######.
                when x"01" & "1100" => d <= "00000000"; -- ........
                when x"01" & "1101" => d <= "00000000"; -- ........
                when x"01" & "1110" => d <= "00000000"; -- ........
                when x"01" & "1111" => d <= "00000000"; -- ........

                when x"02" & "0000" => d <= "00000000"; -- ........
                when x"02" & "0001" => d <= "00000000"; -- ........
                when x"02" & "0010" => d <= "01111110"; -- .######.
                when x"02" & "0011" => d <= "11111111"; -- ########
                when x"02" & "0100" => d <= "11011011"; -- ##.##.##
                when x"02" & "0101" => d <= "11111111"; -- ########
                when x"02" & "0110" => d <= "11111111"; -- ########
                when x"02" & "0111" => d <= "11000011"; -- ##....##
                when x"02" & "1000" => d <= "11100111"; -- ###..###
                when x"02" & "1001" => d <= "11111111"; -- ########
                when x"02" & "1010" => d <= "11111111"; -- ########
                when x"02" & "1011" => d <= "01111110"; -- .######.
                when x"02" & "1100" => d <= "00000000"; -- ........
                when x"02" & "1101" => d <= "00000000"; -- ........
                when x"02" & "1110" => d <= "00000000"; -- ........
                when x"02" & "1111" => d <= "00000000"; -- ........

                when x"03" & "0000" => d <= "00000000"; -- ........
                when x"03" & "0001" => d <= "00000000"; -- ........
                when x"03" & "0010" => d <= "00000000"; -- ........
                when x"03" & "0011" => d <= "00000000"; -- ........
                when x"03" & "0100" => d <= "01101100"; -- .##.##..
                when x"03" & "0101" => d <= "11111110"; -- #######.
                when x"03" & "0110" => d <= "11111110"; -- #######.
                when x"03" & "0111" => d <= "11111110"; -- #######.
                when x"03" & "1000" => d <= "11111110"; -- #######.
                when x"03" & "1001" => d <= "01111100"; -- .#####..
                when x"03" & "1010" => d <= "00111000"; -- ..###...
                when x"03" & "1011" => d <= "00010000"; -- ...#....
                when x"03" & "1100" => d <= "00000000"; -- ........
                when x"03" & "1101" => d <= "00000000"; -- ........
                when x"03" & "1110" => d <= "00000000"; -- ........
                when x"03" & "1111" => d <= "00000000"; -- ........

                when x"04" & "0000" => d <= "00000000"; -- ........
                when x"04" & "0001" => d <= "00000000"; -- ........
                when x"04" & "0010" => d <= "00000000"; -- ........
                when x"04" & "0011" => d <= "00000000"; -- ........
                when x"04" & "0100" => d <= "00010000"; -- ...#....
                when x"04" & "0101" => d <= "00111000"; -- ..###...
                when x"04" & "0110" => d <= "01111100"; -- .#####..
                when x"04" & "0111" => d <= "11111110"; -- #######.
                when x"04" & "1000" => d <= "01111100"; -- .#####..
                when x"04" & "1001" => d <= "00111000"; -- ..###...
                when x"04" & "1010" => d <= "00010000"; -- ...#....
                when x"04" & "1011" => d <= "00000000"; -- ........
                when x"04" & "1100" => d <= "00000000"; -- ........
                when x"04" & "1101" => d <= "00000000"; -- ........
                when x"04" & "1110" => d <= "00000000"; -- ........
                when x"04" & "1111" => d <= "00000000"; -- ........

                when x"05" & "0000" => d <= "00000000"; -- ........
                when x"05" & "0001" => d <= "00000000"; -- ........
                when x"05" & "0010" => d <= "00000000"; -- ........
                when x"05" & "0011" => d <= "00011000"; -- ...##...
                when x"05" & "0100" => d <= "00111100"; -- ..####..
                when x"05" & "0101" => d <= "00111100"; -- ..####..
                when x"05" & "0110" => d <= "11100111"; -- ###..###
                when x"05" & "0111" => d <= "11100111"; -- ###..###
                when x"05" & "1000" => d <= "11100111"; -- ###..###
                when x"05" & "1001" => d <= "00011000"; -- ...##...
                when x"05" & "1010" => d <= "00011000"; -- ...##...
                when x"05" & "1011" => d <= "00111100"; -- ..####..
                when x"05" & "1100" => d <= "00000000"; -- ........
                when x"05" & "1101" => d <= "00000000"; -- ........
                when x"05" & "1110" => d <= "00000000"; -- ........
                when x"05" & "1111" => d <= "00000000"; -- ........

                when x"06" & "0000" => d <= "00000000"; -- ........
                when x"06" & "0001" => d <= "00000000"; -- ........
                when x"06" & "0010" => d <= "00000000"; -- ........
                when x"06" & "0011" => d <= "00011000"; -- ...##...
                when x"06" & "0100" => d <= "00111100"; -- ..####..
                when x"06" & "0101" => d <= "01111110"; -- .######.
                when x"06" & "0110" => d <= "11111111"; -- ########
                when x"06" & "0111" => d <= "11111111"; -- ########
                when x"06" & "1000" => d <= "01111110"; -- .######.
                when x"06" & "1001" => d <= "00011000"; -- ...##...
                when x"06" & "1010" => d <= "00011000"; -- ...##...
                when x"06" & "1011" => d <= "00111100"; -- ..####..
                when x"06" & "1100" => d <= "00000000"; -- ........
                when x"06" & "1101" => d <= "00000000"; -- ........
                when x"06" & "1110" => d <= "00000000"; -- ........
                when x"06" & "1111" => d <= "00000000"; -- ........

                when x"07" & "0000" => d <= "00000000"; -- ........
                when x"07" & "0001" => d <= "00000000"; -- ........
                when x"07" & "0010" => d <= "00000000"; -- ........
                when x"07" & "0011" => d <= "00000000"; -- ........
                when x"07" & "0100" => d <= "00000000"; -- ........
                when x"07" & "0101" => d <= "00000000"; -- ........
                when x"07" & "0110" => d <= "00011000"; -- ...##...
                when x"07" & "0111" => d <= "00111100"; -- ..####..
                when x"07" & "1000" => d <= "00111100"; -- ..####..
                when x"07" & "1001" => d <= "00011000"; -- ...##...
                when x"07" & "1010" => d <= "00000000"; -- ........
                when x"07" & "1011" => d <= "00000000"; -- ........
                when x"07" & "1100" => d <= "00000000"; -- ........
                when x"07" & "1101" => d <= "00000000"; -- ........
                when x"07" & "1110" => d <= "00000000"; -- ........
                when x"07" & "1111" => d <= "00000000"; -- ........

                when x"08" & "0000" => d <= "11111111"; -- ########
                when x"08" & "0001" => d <= "11111111"; -- ########
                when x"08" & "0010" => d <= "11111111"; -- ########
                when x"08" & "0011" => d <= "11111111"; -- ########
                when x"08" & "0100" => d <= "11111111"; -- ########
                when x"08" & "0101" => d <= "11111111"; -- ########
                when x"08" & "0110" => d <= "11100111"; -- ###..###
                when x"08" & "0111" => d <= "11000011"; -- ##....##
                when x"08" & "1000" => d <= "11000011"; -- ##....##
                when x"08" & "1001" => d <= "11100111"; -- ###..###
                when x"08" & "1010" => d <= "11111111"; -- ########
                when x"08" & "1011" => d <= "11111111"; -- ########
                when x"08" & "1100" => d <= "11111111"; -- ########
                when x"08" & "1101" => d <= "11111111"; -- ########
                when x"08" & "1110" => d <= "11111111"; -- ########
                when x"08" & "1111" => d <= "11111111"; -- ########

                when x"09" & "0000" => d <= "00000000"; -- ........
                when x"09" & "0001" => d <= "00000000"; -- ........
                when x"09" & "0010" => d <= "00000000"; -- ........
                when x"09" & "0011" => d <= "00000000"; -- ........
                when x"09" & "0100" => d <= "00000000"; -- ........
                when x"09" & "0101" => d <= "00111100"; -- ..####..
                when x"09" & "0110" => d <= "01100110"; -- .##..##.
                when x"09" & "0111" => d <= "01000010"; -- .#....#.
                when x"09" & "1000" => d <= "01000010"; -- .#....#.
                when x"09" & "1001" => d <= "01100110"; -- .##..##.
                when x"09" & "1010" => d <= "00111100"; -- ..####..
                when x"09" & "1011" => d <= "00000000"; -- ........
                when x"09" & "1100" => d <= "00000000"; -- ........
                when x"09" & "1101" => d <= "00000000"; -- ........
                when x"09" & "1110" => d <= "00000000"; -- ........
                when x"09" & "1111" => d <= "00000000"; -- ........

                when x"0a" & "0000" => d <= "11111111"; -- ########
                when x"0a" & "0001" => d <= "11111111"; -- ########
                when x"0a" & "0010" => d <= "11111111"; -- ########
                when x"0a" & "0011" => d <= "11111111"; -- ########
                when x"0a" & "0100" => d <= "11111111"; -- ########
                when x"0a" & "0101" => d <= "11000011"; -- ##....##
                when x"0a" & "0110" => d <= "10011001"; -- #..##..#
                when x"0a" & "0111" => d <= "10111101"; -- #.####.#
                when x"0a" & "1000" => d <= "10111101"; -- #.####.#
                when x"0a" & "1001" => d <= "10011001"; -- #..##..#
                when x"0a" & "1010" => d <= "11000011"; -- ##....##
                when x"0a" & "1011" => d <= "11111111"; -- ########
                when x"0a" & "1100" => d <= "11111111"; -- ########
                when x"0a" & "1101" => d <= "11111111"; -- ########
                when x"0a" & "1110" => d <= "11111111"; -- ########
                when x"0a" & "1111" => d <= "11111111"; -- ########

                when x"0b" & "0000" => d <= "00000000"; -- ........
                when x"0b" & "0001" => d <= "00000000"; -- ........
                when x"0b" & "0010" => d <= "00011110"; -- ...####.
                when x"0b" & "0011" => d <= "00001110"; -- ....###.
                when x"0b" & "0100" => d <= "00011010"; -- ...##.#.
                when x"0b" & "0101" => d <= "00110010"; -- ..##..#.
                when x"0b" & "0110" => d <= "01111000"; -- .####...
                when x"0b" & "0111" => d <= "11001100"; -- ##..##..
                when x"0b" & "1000" => d <= "11001100"; -- ##..##..
                when x"0b" & "1001" => d <= "11001100"; -- ##..##..
                when x"0b" & "1010" => d <= "11001100"; -- ##..##..
                when x"0b" & "1011" => d <= "01111000"; -- .####...
                when x"0b" & "1100" => d <= "00000000"; -- ........
                when x"0b" & "1101" => d <= "00000000"; -- ........
                when x"0b" & "1110" => d <= "00000000"; -- ........
                when x"0b" & "1111" => d <= "00000000"; -- ........

                when x"0c" & "0000" => d <= "00000000"; -- ........
                when x"0c" & "0001" => d <= "00000000"; -- ........
                when x"0c" & "0010" => d <= "00111100"; -- ..####..
                when x"0c" & "0011" => d <= "01100110"; -- .##..##.
                when x"0c" & "0100" => d <= "01100110"; -- .##..##.
                when x"0c" & "0101" => d <= "01100110"; -- .##..##.
                when x"0c" & "0110" => d <= "01100110"; -- .##..##.
                when x"0c" & "0111" => d <= "00111100"; -- ..####..
                when x"0c" & "1000" => d <= "00011000"; -- ...##...
                when x"0c" & "1001" => d <= "01111110"; -- .######.
                when x"0c" & "1010" => d <= "00011000"; -- ...##...
                when x"0c" & "1011" => d <= "00011000"; -- ...##...
                when x"0c" & "1100" => d <= "00000000"; -- ........
                when x"0c" & "1101" => d <= "00000000"; -- ........
                when x"0c" & "1110" => d <= "00000000"; -- ........
                when x"0c" & "1111" => d <= "00000000"; -- ........

                when x"0d" & "0000" => d <= "00000000"; -- ........
                when x"0d" & "0001" => d <= "00000000"; -- ........
                when x"0d" & "0010" => d <= "00111111"; -- ..######
                when x"0d" & "0011" => d <= "00110011"; -- ..##..##
                when x"0d" & "0100" => d <= "00111111"; -- ..######
                when x"0d" & "0101" => d <= "00110000"; -- ..##....
                when x"0d" & "0110" => d <= "00110000"; -- ..##....
                when x"0d" & "0111" => d <= "00110000"; -- ..##....
                when x"0d" & "1000" => d <= "00110000"; -- ..##....
                when x"0d" & "1001" => d <= "01110000"; -- .###....
                when x"0d" & "1010" => d <= "11110000"; -- ####....
                when x"0d" & "1011" => d <= "11100000"; -- ###.....
                when x"0d" & "1100" => d <= "00000000"; -- ........
                when x"0d" & "1101" => d <= "00000000"; -- ........
                when x"0d" & "1110" => d <= "00000000"; -- ........
                when x"0d" & "1111" => d <= "00000000"; -- ........

                when x"0e" & "0000" => d <= "00000000"; -- ........
                when x"0e" & "0001" => d <= "00000000"; -- ........
                when x"0e" & "0010" => d <= "01111111"; -- .#######
                when x"0e" & "0011" => d <= "01100011"; -- .##...##
                when x"0e" & "0100" => d <= "01111111"; -- .#######
                when x"0e" & "0101" => d <= "01100011"; -- .##...##
                when x"0e" & "0110" => d <= "01100011"; -- .##...##
                when x"0e" & "0111" => d <= "01100011"; -- .##...##
                when x"0e" & "1000" => d <= "01100011"; -- .##...##
                when x"0e" & "1001" => d <= "01100111"; -- .##..###
                when x"0e" & "1010" => d <= "11100111"; -- ###..###
                when x"0e" & "1011" => d <= "11100110"; -- ###..##.
                when x"0e" & "1100" => d <= "11000000"; -- ##......
                when x"0e" & "1101" => d <= "00000000"; -- ........
                when x"0e" & "1110" => d <= "00000000"; -- ........
                when x"0e" & "1111" => d <= "00000000"; -- ........

                when x"0f" & "0000" => d <= "00000000"; -- ........
                when x"0f" & "0001" => d <= "00000000"; -- ........
                when x"0f" & "0010" => d <= "00000000"; -- ........
                when x"0f" & "0011" => d <= "00011000"; -- ...##...
                when x"0f" & "0100" => d <= "00011000"; -- ...##...
                when x"0f" & "0101" => d <= "11011011"; -- ##.##.##
                when x"0f" & "0110" => d <= "00111100"; -- ..####..
                when x"0f" & "0111" => d <= "11100111"; -- ###..###
                when x"0f" & "1000" => d <= "00111100"; -- ..####..
                when x"0f" & "1001" => d <= "11011011"; -- ##.##.##
                when x"0f" & "1010" => d <= "00011000"; -- ...##...
                when x"0f" & "1011" => d <= "00011000"; -- ...##...
                when x"0f" & "1100" => d <= "00000000"; -- ........
                when x"0f" & "1101" => d <= "00000000"; -- ........
                when x"0f" & "1110" => d <= "00000000"; -- ........
                when x"0f" & "1111" => d <= "00000000"; -- ........

                when x"10" & "0000" => d <= "00000000"; -- ........
                when x"10" & "0001" => d <= "10000000"; -- #.......
                when x"10" & "0010" => d <= "11000000"; -- ##......
                when x"10" & "0011" => d <= "11100000"; -- ###.....
                when x"10" & "0100" => d <= "11110000"; -- ####....
                when x"10" & "0101" => d <= "11111000"; -- #####...
                when x"10" & "0110" => d <= "11111110"; -- #######.
                when x"10" & "0111" => d <= "11111000"; -- #####...
                when x"10" & "1000" => d <= "11110000"; -- ####....
                when x"10" & "1001" => d <= "11100000"; -- ###.....
                when x"10" & "1010" => d <= "11000000"; -- ##......
                when x"10" & "1011" => d <= "10000000"; -- #.......
                when x"10" & "1100" => d <= "00000000"; -- ........
                when x"10" & "1101" => d <= "00000000"; -- ........
                when x"10" & "1110" => d <= "00000000"; -- ........
                when x"10" & "1111" => d <= "00000000"; -- ........

                when x"11" & "0000" => d <= "00000000"; -- ........
                when x"11" & "0001" => d <= "00000010"; -- ......#.
                when x"11" & "0010" => d <= "00000110"; -- .....##.
                when x"11" & "0011" => d <= "00001110"; -- ....###.
                when x"11" & "0100" => d <= "00011110"; -- ...####.
                when x"11" & "0101" => d <= "00111110"; -- ..#####.
                when x"11" & "0110" => d <= "11111110"; -- #######.
                when x"11" & "0111" => d <= "00111110"; -- ..#####.
                when x"11" & "1000" => d <= "00011110"; -- ...####.
                when x"11" & "1001" => d <= "00001110"; -- ....###.
                when x"11" & "1010" => d <= "00000110"; -- .....##.
                when x"11" & "1011" => d <= "00000010"; -- ......#.
                when x"11" & "1100" => d <= "00000000"; -- ........
                when x"11" & "1101" => d <= "00000000"; -- ........
                when x"11" & "1110" => d <= "00000000"; -- ........
                when x"11" & "1111" => d <= "00000000"; -- ........

                when x"12" & "0000" => d <= "00000000"; -- ........
                when x"12" & "0001" => d <= "00000000"; -- ........
                when x"12" & "0010" => d <= "00011000"; -- ...##...
                when x"12" & "0011" => d <= "00111100"; -- ..####..
                when x"12" & "0100" => d <= "01111110"; -- .######.
                when x"12" & "0101" => d <= "00011000"; -- ...##...
                when x"12" & "0110" => d <= "00011000"; -- ...##...
                when x"12" & "0111" => d <= "00011000"; -- ...##...
                when x"12" & "1000" => d <= "01111110"; -- .######.
                when x"12" & "1001" => d <= "00111100"; -- ..####..
                when x"12" & "1010" => d <= "00011000"; -- ...##...
                when x"12" & "1011" => d <= "00000000"; -- ........
                when x"12" & "1100" => d <= "00000000"; -- ........
                when x"12" & "1101" => d <= "00000000"; -- ........
                when x"12" & "1110" => d <= "00000000"; -- ........
                when x"12" & "1111" => d <= "00000000"; -- ........

                when x"13" & "0000" => d <= "00000000"; -- ........
                when x"13" & "0001" => d <= "00000000"; -- ........
                when x"13" & "0010" => d <= "01100110"; -- .##..##.
                when x"13" & "0011" => d <= "01100110"; -- .##..##.
                when x"13" & "0100" => d <= "01100110"; -- .##..##.
                when x"13" & "0101" => d <= "01100110"; -- .##..##.
                when x"13" & "0110" => d <= "01100110"; -- .##..##.
                when x"13" & "0111" => d <= "01100110"; -- .##..##.
                when x"13" & "1000" => d <= "01100110"; -- .##..##.
                when x"13" & "1001" => d <= "00000000"; -- ........
                when x"13" & "1010" => d <= "01100110"; -- .##..##.
                when x"13" & "1011" => d <= "01100110"; -- .##..##.
                when x"13" & "1100" => d <= "00000000"; -- ........
                when x"13" & "1101" => d <= "00000000"; -- ........
                when x"13" & "1110" => d <= "00000000"; -- ........
                when x"13" & "1111" => d <= "00000000"; -- ........

                when x"14" & "0000" => d <= "00000000"; -- ........
                when x"14" & "0001" => d <= "00000000"; -- ........
                when x"14" & "0010" => d <= "01111111"; -- .#######
                when x"14" & "0011" => d <= "11011011"; -- ##.##.##
                when x"14" & "0100" => d <= "11011011"; -- ##.##.##
                when x"14" & "0101" => d <= "11011011"; -- ##.##.##
                when x"14" & "0110" => d <= "01111011"; -- .####.##
                when x"14" & "0111" => d <= "00011011"; -- ...##.##
                when x"14" & "1000" => d <= "00011011"; -- ...##.##
                when x"14" & "1001" => d <= "00011011"; -- ...##.##
                when x"14" & "1010" => d <= "00011011"; -- ...##.##
                when x"14" & "1011" => d <= "00011011"; -- ...##.##
                when x"14" & "1100" => d <= "00000000"; -- ........
                when x"14" & "1101" => d <= "00000000"; -- ........
                when x"14" & "1110" => d <= "00000000"; -- ........
                when x"14" & "1111" => d <= "00000000"; -- ........

                when x"15" & "0000" => d <= "00000000"; -- ........
                when x"15" & "0001" => d <= "01111100"; -- .#####..
                when x"15" & "0010" => d <= "11000110"; -- ##...##.
                when x"15" & "0011" => d <= "01100000"; -- .##.....
                when x"15" & "0100" => d <= "00111000"; -- ..###...
                when x"15" & "0101" => d <= "01101100"; -- .##.##..
                when x"15" & "0110" => d <= "11000110"; -- ##...##.
                when x"15" & "0111" => d <= "11000110"; -- ##...##.
                when x"15" & "1000" => d <= "01101100"; -- .##.##..
                when x"15" & "1001" => d <= "00111000"; -- ..###...
                when x"15" & "1010" => d <= "00001100"; -- ....##..
                when x"15" & "1011" => d <= "11000110"; -- ##...##.
                when x"15" & "1100" => d <= "01111100"; -- .#####..
                when x"15" & "1101" => d <= "00000000"; -- ........
                when x"15" & "1110" => d <= "00000000"; -- ........
                when x"15" & "1111" => d <= "00000000"; -- ........

                when x"16" & "0000" => d <= "00000000"; -- ........
                when x"16" & "0001" => d <= "00000000"; -- ........
                when x"16" & "0010" => d <= "00000000"; -- ........
                when x"16" & "0011" => d <= "00000000"; -- ........
                when x"16" & "0100" => d <= "00000000"; -- ........
                when x"16" & "0101" => d <= "00000000"; -- ........
                when x"16" & "0110" => d <= "00000000"; -- ........
                when x"16" & "0111" => d <= "00000000"; -- ........
                when x"16" & "1000" => d <= "11111110"; -- #######.
                when x"16" & "1001" => d <= "11111110"; -- #######.
                when x"16" & "1010" => d <= "11111110"; -- #######.
                when x"16" & "1011" => d <= "11111110"; -- #######.
                when x"16" & "1100" => d <= "00000000"; -- ........
                when x"16" & "1101" => d <= "00000000"; -- ........
                when x"16" & "1110" => d <= "00000000"; -- ........
                when x"16" & "1111" => d <= "00000000"; -- ........

                when x"17" & "0000" => d <= "00000000"; -- ........
                when x"17" & "0001" => d <= "00000000"; -- ........
                when x"17" & "0010" => d <= "00011000"; -- ...##...
                when x"17" & "0011" => d <= "00111100"; -- ..####..
                when x"17" & "0100" => d <= "01111110"; -- .######.
                when x"17" & "0101" => d <= "00011000"; -- ...##...
                when x"17" & "0110" => d <= "00011000"; -- ...##...
                when x"17" & "0111" => d <= "00011000"; -- ...##...
                when x"17" & "1000" => d <= "01111110"; -- .######.
                when x"17" & "1001" => d <= "00111100"; -- ..####..
                when x"17" & "1010" => d <= "00011000"; -- ...##...
                when x"17" & "1011" => d <= "01111110"; -- .######.
                when x"17" & "1100" => d <= "00000000"; -- ........
                when x"17" & "1101" => d <= "00000000"; -- ........
                when x"17" & "1110" => d <= "00000000"; -- ........
                when x"17" & "1111" => d <= "00000000"; -- ........

                when x"18" & "0000" => d <= "00000000"; -- ........
                when x"18" & "0001" => d <= "00000000"; -- ........
                when x"18" & "0010" => d <= "00011000"; -- ...##...
                when x"18" & "0011" => d <= "00111100"; -- ..####..
                when x"18" & "0100" => d <= "01111110"; -- .######.
                when x"18" & "0101" => d <= "00011000"; -- ...##...
                when x"18" & "0110" => d <= "00011000"; -- ...##...
                when x"18" & "0111" => d <= "00011000"; -- ...##...
                when x"18" & "1000" => d <= "00011000"; -- ...##...
                when x"18" & "1001" => d <= "00011000"; -- ...##...
                when x"18" & "1010" => d <= "00011000"; -- ...##...
                when x"18" & "1011" => d <= "00011000"; -- ...##...
                when x"18" & "1100" => d <= "00000000"; -- ........
                when x"18" & "1101" => d <= "00000000"; -- ........
                when x"18" & "1110" => d <= "00000000"; -- ........
                when x"18" & "1111" => d <= "00000000"; -- ........

                when x"19" & "0000" => d <= "00000000"; -- ........
                when x"19" & "0001" => d <= "00000000"; -- ........
                when x"19" & "0010" => d <= "00011000"; -- ...##...
                when x"19" & "0011" => d <= "00011000"; -- ...##...
                when x"19" & "0100" => d <= "00011000"; -- ...##...
                when x"19" & "0101" => d <= "00011000"; -- ...##...
                when x"19" & "0110" => d <= "00011000"; -- ...##...
                when x"19" & "0111" => d <= "00011000"; -- ...##...
                when x"19" & "1000" => d <= "00011000"; -- ...##...
                when x"19" & "1001" => d <= "01111110"; -- .######.
                when x"19" & "1010" => d <= "00111100"; -- ..####..
                when x"19" & "1011" => d <= "00011000"; -- ...##...
                when x"19" & "1100" => d <= "00000000"; -- ........
                when x"19" & "1101" => d <= "00000000"; -- ........
                when x"19" & "1110" => d <= "00000000"; -- ........
                when x"19" & "1111" => d <= "00000000"; -- ........

                when x"1a" & "0000" => d <= "00000000"; -- ........
                when x"1a" & "0001" => d <= "00000000"; -- ........
                when x"1a" & "0010" => d <= "00000000"; -- ........
                when x"1a" & "0011" => d <= "00000000"; -- ........
                when x"1a" & "0100" => d <= "00000000"; -- ........
                when x"1a" & "0101" => d <= "00011000"; -- ...##...
                when x"1a" & "0110" => d <= "00001100"; -- ....##..
                when x"1a" & "0111" => d <= "11111110"; -- #######.
                when x"1a" & "1000" => d <= "00001100"; -- ....##..
                when x"1a" & "1001" => d <= "00011000"; -- ...##...
                when x"1a" & "1010" => d <= "00000000"; -- ........
                when x"1a" & "1011" => d <= "00000000"; -- ........
                when x"1a" & "1100" => d <= "00000000"; -- ........
                when x"1a" & "1101" => d <= "00000000"; -- ........
                when x"1a" & "1110" => d <= "00000000"; -- ........
                when x"1a" & "1111" => d <= "00000000"; -- ........

                when x"1b" & "0000" => d <= "00000000"; -- ........
                when x"1b" & "0001" => d <= "00000000"; -- ........
                when x"1b" & "0010" => d <= "00000000"; -- ........
                when x"1b" & "0011" => d <= "00000000"; -- ........
                when x"1b" & "0100" => d <= "00000000"; -- ........
                when x"1b" & "0101" => d <= "00110000"; -- ..##....
                when x"1b" & "0110" => d <= "01100000"; -- .##.....
                when x"1b" & "0111" => d <= "11111110"; -- #######.
                when x"1b" & "1000" => d <= "01100000"; -- .##.....
                when x"1b" & "1001" => d <= "00110000"; -- ..##....
                when x"1b" & "1010" => d <= "00000000"; -- ........
                when x"1b" & "1011" => d <= "00000000"; -- ........
                when x"1b" & "1100" => d <= "00000000"; -- ........
                when x"1b" & "1101" => d <= "00000000"; -- ........
                when x"1b" & "1110" => d <= "00000000"; -- ........
                when x"1b" & "1111" => d <= "00000000"; -- ........

                when x"1c" & "0000" => d <= "00000000"; -- ........
                when x"1c" & "0001" => d <= "00000000"; -- ........
                when x"1c" & "0010" => d <= "00000000"; -- ........
                when x"1c" & "0011" => d <= "00000000"; -- ........
                when x"1c" & "0100" => d <= "00000000"; -- ........
                when x"1c" & "0101" => d <= "00000000"; -- ........
                when x"1c" & "0110" => d <= "11000000"; -- ##......
                when x"1c" & "0111" => d <= "11000000"; -- ##......
                when x"1c" & "1000" => d <= "11000000"; -- ##......
                when x"1c" & "1001" => d <= "11111110"; -- #######.
                when x"1c" & "1010" => d <= "00000000"; -- ........
                when x"1c" & "1011" => d <= "00000000"; -- ........
                when x"1c" & "1100" => d <= "00000000"; -- ........
                when x"1c" & "1101" => d <= "00000000"; -- ........
                when x"1c" & "1110" => d <= "00000000"; -- ........
                when x"1c" & "1111" => d <= "00000000"; -- ........

                when x"1d" & "0000" => d <= "00000000"; -- ........
                when x"1d" & "0001" => d <= "00000000"; -- ........
                when x"1d" & "0010" => d <= "00000000"; -- ........
                when x"1d" & "0011" => d <= "00000000"; -- ........
                when x"1d" & "0100" => d <= "00000000"; -- ........
                when x"1d" & "0101" => d <= "00101000"; -- ..#.#...
                when x"1d" & "0110" => d <= "01101100"; -- .##.##..
                when x"1d" & "0111" => d <= "11111110"; -- #######.
                when x"1d" & "1000" => d <= "01101100"; -- .##.##..
                when x"1d" & "1001" => d <= "00101000"; -- ..#.#...
                when x"1d" & "1010" => d <= "00000000"; -- ........
                when x"1d" & "1011" => d <= "00000000"; -- ........
                when x"1d" & "1100" => d <= "00000000"; -- ........
                when x"1d" & "1101" => d <= "00000000"; -- ........
                when x"1d" & "1110" => d <= "00000000"; -- ........
                when x"1d" & "1111" => d <= "00000000"; -- ........

                when x"1e" & "0000" => d <= "00000000"; -- ........
                when x"1e" & "0001" => d <= "00000000"; -- ........
                when x"1e" & "0010" => d <= "00000000"; -- ........
                when x"1e" & "0011" => d <= "00000000"; -- ........
                when x"1e" & "0100" => d <= "00010000"; -- ...#....
                when x"1e" & "0101" => d <= "00111000"; -- ..###...
                when x"1e" & "0110" => d <= "00111000"; -- ..###...
                when x"1e" & "0111" => d <= "01111100"; -- .#####..
                when x"1e" & "1000" => d <= "01111100"; -- .#####..
                when x"1e" & "1001" => d <= "11111110"; -- #######.
                when x"1e" & "1010" => d <= "11111110"; -- #######.
                when x"1e" & "1011" => d <= "00000000"; -- ........
                when x"1e" & "1100" => d <= "00000000"; -- ........
                when x"1e" & "1101" => d <= "00000000"; -- ........
                when x"1e" & "1110" => d <= "00000000"; -- ........
                when x"1e" & "1111" => d <= "00000000"; -- ........

                when x"1f" & "0000" => d <= "00000000"; -- ........
                when x"1f" & "0001" => d <= "00000000"; -- ........
                when x"1f" & "0010" => d <= "00000000"; -- ........
                when x"1f" & "0011" => d <= "00000000"; -- ........
                when x"1f" & "0100" => d <= "11111110"; -- #######.
                when x"1f" & "0101" => d <= "11111110"; -- #######.
                when x"1f" & "0110" => d <= "01111100"; -- .#####..
                when x"1f" & "0111" => d <= "01111100"; -- .#####..
                when x"1f" & "1000" => d <= "00111000"; -- ..###...
                when x"1f" & "1001" => d <= "00111000"; -- ..###...
                when x"1f" & "1010" => d <= "00010000"; -- ...#....
                when x"1f" & "1011" => d <= "00000000"; -- ........
                when x"1f" & "1100" => d <= "00000000"; -- ........
                when x"1f" & "1101" => d <= "00000000"; -- ........
                when x"1f" & "1110" => d <= "00000000"; -- ........
                when x"1f" & "1111" => d <= "00000000"; -- ........

                when x"20" & "0000" => d <= "00000000"; -- ........
                when x"20" & "0001" => d <= "00000000"; -- ........
                when x"20" & "0010" => d <= "00000000"; -- ........
                when x"20" & "0011" => d <= "00000000"; -- ........
                when x"20" & "0100" => d <= "00000000"; -- ........
                when x"20" & "0101" => d <= "00000000"; -- ........
                when x"20" & "0110" => d <= "00000000"; -- ........
                when x"20" & "0111" => d <= "00000000"; -- ........
                when x"20" & "1000" => d <= "00000000"; -- ........
                when x"20" & "1001" => d <= "00000000"; -- ........
                when x"20" & "1010" => d <= "00000000"; -- ........
                when x"20" & "1011" => d <= "00000000"; -- ........
                when x"20" & "1100" => d <= "00000000"; -- ........
                when x"20" & "1101" => d <= "00000000"; -- ........
                when x"20" & "1110" => d <= "00000000"; -- ........
                when x"20" & "1111" => d <= "00000000"; -- ........

                when x"21" & "0000" => d <= "00000000"; -- ........
                when x"21" & "0001" => d <= "00000000"; -- ........
                when x"21" & "0010" => d <= "00011000"; -- ...##...
                when x"21" & "0011" => d <= "00111100"; -- ..####..
                when x"21" & "0100" => d <= "00111100"; -- ..####..
                when x"21" & "0101" => d <= "00111100"; -- ..####..
                when x"21" & "0110" => d <= "00011000"; -- ...##...
                when x"21" & "0111" => d <= "00011000"; -- ...##...
                when x"21" & "1000" => d <= "00011000"; -- ...##...
                when x"21" & "1001" => d <= "00000000"; -- ........
                when x"21" & "1010" => d <= "00011000"; -- ...##...
                when x"21" & "1011" => d <= "00011000"; -- ...##...
                when x"21" & "1100" => d <= "00000000"; -- ........
                when x"21" & "1101" => d <= "00000000"; -- ........
                when x"21" & "1110" => d <= "00000000"; -- ........
                when x"21" & "1111" => d <= "00000000"; -- ........

                when x"22" & "0000" => d <= "00000000"; -- ........
                when x"22" & "0001" => d <= "01100110"; -- .##..##.
                when x"22" & "0010" => d <= "01100110"; -- .##..##.
                when x"22" & "0011" => d <= "01100110"; -- .##..##.
                when x"22" & "0100" => d <= "00100100"; -- ..#..#..
                when x"22" & "0101" => d <= "00000000"; -- ........
                when x"22" & "0110" => d <= "00000000"; -- ........
                when x"22" & "0111" => d <= "00000000"; -- ........
                when x"22" & "1000" => d <= "00000000"; -- ........
                when x"22" & "1001" => d <= "00000000"; -- ........
                when x"22" & "1010" => d <= "00000000"; -- ........
                when x"22" & "1011" => d <= "00000000"; -- ........
                when x"22" & "1100" => d <= "00000000"; -- ........
                when x"22" & "1101" => d <= "00000000"; -- ........
                when x"22" & "1110" => d <= "00000000"; -- ........
                when x"22" & "1111" => d <= "00000000"; -- ........

                when x"23" & "0000" => d <= "00000000"; -- ........
                when x"23" & "0001" => d <= "00000000"; -- ........
                when x"23" & "0010" => d <= "00000000"; -- ........
                when x"23" & "0011" => d <= "01101100"; -- .##.##..
                when x"23" & "0100" => d <= "01101100"; -- .##.##..
                when x"23" & "0101" => d <= "11111110"; -- #######.
                when x"23" & "0110" => d <= "01101100"; -- .##.##..
                when x"23" & "0111" => d <= "01101100"; -- .##.##..
                when x"23" & "1000" => d <= "01101100"; -- .##.##..
                when x"23" & "1001" => d <= "11111110"; -- #######.
                when x"23" & "1010" => d <= "01101100"; -- .##.##..
                when x"23" & "1011" => d <= "01101100"; -- .##.##..
                when x"23" & "1100" => d <= "00000000"; -- ........
                when x"23" & "1101" => d <= "00000000"; -- ........
                when x"23" & "1110" => d <= "00000000"; -- ........
                when x"23" & "1111" => d <= "00000000"; -- ........

                when x"24" & "0000" => d <= "00011000"; -- ...##...
                when x"24" & "0001" => d <= "00011000"; -- ...##...
                when x"24" & "0010" => d <= "01111100"; -- .#####..
                when x"24" & "0011" => d <= "11000110"; -- ##...##.
                when x"24" & "0100" => d <= "11000010"; -- ##....#.
                when x"24" & "0101" => d <= "11000000"; -- ##......
                when x"24" & "0110" => d <= "01111100"; -- .#####..
                when x"24" & "0111" => d <= "00000110"; -- .....##.
                when x"24" & "1000" => d <= "00000110"; -- .....##.
                when x"24" & "1001" => d <= "10000110"; -- #....##.
                when x"24" & "1010" => d <= "11000110"; -- ##...##.
                when x"24" & "1011" => d <= "01111100"; -- .#####..
                when x"24" & "1100" => d <= "00011000"; -- ...##...
                when x"24" & "1101" => d <= "00011000"; -- ...##...
                when x"24" & "1110" => d <= "00000000"; -- ........
                when x"24" & "1111" => d <= "00000000"; -- ........

                when x"25" & "0000" => d <= "00000000"; -- ........
                when x"25" & "0001" => d <= "00000000"; -- ........
                when x"25" & "0010" => d <= "00000000"; -- ........
                when x"25" & "0011" => d <= "00000000"; -- ........
                when x"25" & "0100" => d <= "11000010"; -- ##....#.
                when x"25" & "0101" => d <= "11000110"; -- ##...##.
                when x"25" & "0110" => d <= "00001100"; -- ....##..
                when x"25" & "0111" => d <= "00011000"; -- ...##...
                when x"25" & "1000" => d <= "00110000"; -- ..##....
                when x"25" & "1001" => d <= "01100000"; -- .##.....
                when x"25" & "1010" => d <= "11000110"; -- ##...##.
                when x"25" & "1011" => d <= "10000110"; -- #....##.
                when x"25" & "1100" => d <= "00000000"; -- ........
                when x"25" & "1101" => d <= "00000000"; -- ........
                when x"25" & "1110" => d <= "00000000"; -- ........
                when x"25" & "1111" => d <= "00000000"; -- ........

                when x"26" & "0000" => d <= "00000000"; -- ........
                when x"26" & "0001" => d <= "00000000"; -- ........
                when x"26" & "0010" => d <= "00111000"; -- ..###...
                when x"26" & "0011" => d <= "01101100"; -- .##.##..
                when x"26" & "0100" => d <= "01101100"; -- .##.##..
                when x"26" & "0101" => d <= "00111000"; -- ..###...
                when x"26" & "0110" => d <= "01110110"; -- .###.##.
                when x"26" & "0111" => d <= "11011100"; -- ##.###..
                when x"26" & "1000" => d <= "11001100"; -- ##..##..
                when x"26" & "1001" => d <= "11001100"; -- ##..##..
                when x"26" & "1010" => d <= "11001100"; -- ##..##..
                when x"26" & "1011" => d <= "01110110"; -- .###.##.
                when x"26" & "1100" => d <= "00000000"; -- ........
                when x"26" & "1101" => d <= "00000000"; -- ........
                when x"26" & "1110" => d <= "00000000"; -- ........
                when x"26" & "1111" => d <= "00000000"; -- ........

                when x"27" & "0000" => d <= "00000000"; -- ........
                when x"27" & "0001" => d <= "00110000"; -- ..##....
                when x"27" & "0010" => d <= "00110000"; -- ..##....
                when x"27" & "0011" => d <= "00110000"; -- ..##....
                when x"27" & "0100" => d <= "01100000"; -- .##.....
                when x"27" & "0101" => d <= "00000000"; -- ........
                when x"27" & "0110" => d <= "00000000"; -- ........
                when x"27" & "0111" => d <= "00000000"; -- ........
                when x"27" & "1000" => d <= "00000000"; -- ........
                when x"27" & "1001" => d <= "00000000"; -- ........
                when x"27" & "1010" => d <= "00000000"; -- ........
                when x"27" & "1011" => d <= "00000000"; -- ........
                when x"27" & "1100" => d <= "00000000"; -- ........
                when x"27" & "1101" => d <= "00000000"; -- ........
                when x"27" & "1110" => d <= "00000000"; -- ........
                when x"27" & "1111" => d <= "00000000"; -- ........

                when x"28" & "0000" => d <= "00000000"; -- ........
                when x"28" & "0001" => d <= "00000000"; -- ........
                when x"28" & "0010" => d <= "00001100"; -- ....##..
                when x"28" & "0011" => d <= "00011000"; -- ...##...
                when x"28" & "0100" => d <= "00110000"; -- ..##....
                when x"28" & "0101" => d <= "00110000"; -- ..##....
                when x"28" & "0110" => d <= "00110000"; -- ..##....
                when x"28" & "0111" => d <= "00110000"; -- ..##....
                when x"28" & "1000" => d <= "00110000"; -- ..##....
                when x"28" & "1001" => d <= "00110000"; -- ..##....
                when x"28" & "1010" => d <= "00011000"; -- ...##...
                when x"28" & "1011" => d <= "00001100"; -- ....##..
                when x"28" & "1100" => d <= "00000000"; -- ........
                when x"28" & "1101" => d <= "00000000"; -- ........
                when x"28" & "1110" => d <= "00000000"; -- ........
                when x"28" & "1111" => d <= "00000000"; -- ........

                when x"29" & "0000" => d <= "00000000"; -- ........
                when x"29" & "0001" => d <= "00000000"; -- ........
                when x"29" & "0010" => d <= "00110000"; -- ..##....
                when x"29" & "0011" => d <= "00011000"; -- ...##...
                when x"29" & "0100" => d <= "00001100"; -- ....##..
                when x"29" & "0101" => d <= "00001100"; -- ....##..
                when x"29" & "0110" => d <= "00001100"; -- ....##..
                when x"29" & "0111" => d <= "00001100"; -- ....##..
                when x"29" & "1000" => d <= "00001100"; -- ....##..
                when x"29" & "1001" => d <= "00001100"; -- ....##..
                when x"29" & "1010" => d <= "00011000"; -- ...##...
                when x"29" & "1011" => d <= "00110000"; -- ..##....
                when x"29" & "1100" => d <= "00000000"; -- ........
                when x"29" & "1101" => d <= "00000000"; -- ........
                when x"29" & "1110" => d <= "00000000"; -- ........
                when x"29" & "1111" => d <= "00000000"; -- ........

                when x"2a" & "0000" => d <= "00000000"; -- ........
                when x"2a" & "0001" => d <= "00000000"; -- ........
                when x"2a" & "0010" => d <= "00000000"; -- ........
                when x"2a" & "0011" => d <= "00000000"; -- ........
                when x"2a" & "0100" => d <= "00000000"; -- ........
                when x"2a" & "0101" => d <= "01100110"; -- .##..##.
                when x"2a" & "0110" => d <= "00111100"; -- ..####..
                when x"2a" & "0111" => d <= "11111111"; -- ########
                when x"2a" & "1000" => d <= "00111100"; -- ..####..
                when x"2a" & "1001" => d <= "01100110"; -- .##..##.
                when x"2a" & "1010" => d <= "00000000"; -- ........
                when x"2a" & "1011" => d <= "00000000"; -- ........
                when x"2a" & "1100" => d <= "00000000"; -- ........
                when x"2a" & "1101" => d <= "00000000"; -- ........
                when x"2a" & "1110" => d <= "00000000"; -- ........
                when x"2a" & "1111" => d <= "00000000"; -- ........

                when x"2b" & "0000" => d <= "00000000"; -- ........
                when x"2b" & "0001" => d <= "00000000"; -- ........
                when x"2b" & "0010" => d <= "00000000"; -- ........
                when x"2b" & "0011" => d <= "00000000"; -- ........
                when x"2b" & "0100" => d <= "00000000"; -- ........
                when x"2b" & "0101" => d <= "00011000"; -- ...##...
                when x"2b" & "0110" => d <= "00011000"; -- ...##...
                when x"2b" & "0111" => d <= "01111110"; -- .######.
                when x"2b" & "1000" => d <= "00011000"; -- ...##...
                when x"2b" & "1001" => d <= "00011000"; -- ...##...
                when x"2b" & "1010" => d <= "00000000"; -- ........
                when x"2b" & "1011" => d <= "00000000"; -- ........
                when x"2b" & "1100" => d <= "00000000"; -- ........
                when x"2b" & "1101" => d <= "00000000"; -- ........
                when x"2b" & "1110" => d <= "00000000"; -- ........
                when x"2b" & "1111" => d <= "00000000"; -- ........

                when x"2c" & "0000" => d <= "00000000"; -- ........
                when x"2c" & "0001" => d <= "00000000"; -- ........
                when x"2c" & "0010" => d <= "00000000"; -- ........
                when x"2c" & "0011" => d <= "00000000"; -- ........
                when x"2c" & "0100" => d <= "00000000"; -- ........
                when x"2c" & "0101" => d <= "00000000"; -- ........
                when x"2c" & "0110" => d <= "00000000"; -- ........
                when x"2c" & "0111" => d <= "00000000"; -- ........
                when x"2c" & "1000" => d <= "00000000"; -- ........
                when x"2c" & "1001" => d <= "00011000"; -- ...##...
                when x"2c" & "1010" => d <= "00011000"; -- ...##...
                when x"2c" & "1011" => d <= "00011000"; -- ...##...
                when x"2c" & "1100" => d <= "00110000"; -- ..##....
                when x"2c" & "1101" => d <= "00000000"; -- ........
                when x"2c" & "1110" => d <= "00000000"; -- ........
                when x"2c" & "1111" => d <= "00000000"; -- ........

                when x"2d" & "0000" => d <= "00000000"; -- ........
                when x"2d" & "0001" => d <= "00000000"; -- ........
                when x"2d" & "0010" => d <= "00000000"; -- ........
                when x"2d" & "0011" => d <= "00000000"; -- ........
                when x"2d" & "0100" => d <= "00000000"; -- ........
                when x"2d" & "0101" => d <= "00000000"; -- ........
                when x"2d" & "0110" => d <= "00000000"; -- ........
                when x"2d" & "0111" => d <= "11111110"; -- #######.
                when x"2d" & "1000" => d <= "00000000"; -- ........
                when x"2d" & "1001" => d <= "00000000"; -- ........
                when x"2d" & "1010" => d <= "00000000"; -- ........
                when x"2d" & "1011" => d <= "00000000"; -- ........
                when x"2d" & "1100" => d <= "00000000"; -- ........
                when x"2d" & "1101" => d <= "00000000"; -- ........
                when x"2d" & "1110" => d <= "00000000"; -- ........
                when x"2d" & "1111" => d <= "00000000"; -- ........

                when x"2e" & "0000" => d <= "00000000"; -- ........
                when x"2e" & "0001" => d <= "00000000"; -- ........
                when x"2e" & "0010" => d <= "00000000"; -- ........
                when x"2e" & "0011" => d <= "00000000"; -- ........
                when x"2e" & "0100" => d <= "00000000"; -- ........
                when x"2e" & "0101" => d <= "00000000"; -- ........
                when x"2e" & "0110" => d <= "00000000"; -- ........
                when x"2e" & "0111" => d <= "00000000"; -- ........
                when x"2e" & "1000" => d <= "00000000"; -- ........
                when x"2e" & "1001" => d <= "00000000"; -- ........
                when x"2e" & "1010" => d <= "00011000"; -- ...##...
                when x"2e" & "1011" => d <= "00011000"; -- ...##...
                when x"2e" & "1100" => d <= "00000000"; -- ........
                when x"2e" & "1101" => d <= "00000000"; -- ........
                when x"2e" & "1110" => d <= "00000000"; -- ........
                when x"2e" & "1111" => d <= "00000000"; -- ........

                when x"2f" & "0000" => d <= "00000000"; -- ........
                when x"2f" & "0001" => d <= "00000000"; -- ........
                when x"2f" & "0010" => d <= "00000000"; -- ........
                when x"2f" & "0011" => d <= "00000000"; -- ........
                when x"2f" & "0100" => d <= "00000010"; -- ......#.
                when x"2f" & "0101" => d <= "00000110"; -- .....##.
                when x"2f" & "0110" => d <= "00001100"; -- ....##..
                when x"2f" & "0111" => d <= "00011000"; -- ...##...
                when x"2f" & "1000" => d <= "00110000"; -- ..##....
                when x"2f" & "1001" => d <= "01100000"; -- .##.....
                when x"2f" & "1010" => d <= "11000000"; -- ##......
                when x"2f" & "1011" => d <= "10000000"; -- #.......
                when x"2f" & "1100" => d <= "00000000"; -- ........
                when x"2f" & "1101" => d <= "00000000"; -- ........
                when x"2f" & "1110" => d <= "00000000"; -- ........
                when x"2f" & "1111" => d <= "00000000"; -- ........

                when x"30" & "0000" => d <= "00000000"; -- ........
                when x"30" & "0001" => d <= "00000000"; -- ........
                when x"30" & "0010" => d <= "00111000"; -- ..###...
                when x"30" & "0011" => d <= "01101100"; -- .##.##..
                when x"30" & "0100" => d <= "11000110"; -- ##...##.
                when x"30" & "0101" => d <= "11000110"; -- ##...##.
                when x"30" & "0110" => d <= "11010110"; -- ##.#.##.
                when x"30" & "0111" => d <= "11010110"; -- ##.#.##.
                when x"30" & "1000" => d <= "11000110"; -- ##...##.
                when x"30" & "1001" => d <= "11000110"; -- ##...##.
                when x"30" & "1010" => d <= "01101100"; -- .##.##..
                when x"30" & "1011" => d <= "00111000"; -- ..###...
                when x"30" & "1100" => d <= "00000000"; -- ........
                when x"30" & "1101" => d <= "00000000"; -- ........
                when x"30" & "1110" => d <= "00000000"; -- ........
                when x"30" & "1111" => d <= "00000000"; -- ........

                when x"31" & "0000" => d <= "00000000"; -- ........
                when x"31" & "0001" => d <= "00000000"; -- ........
                when x"31" & "0010" => d <= "00011000"; -- ...##...
                when x"31" & "0011" => d <= "00111000"; -- ..###...
                when x"31" & "0100" => d <= "01111000"; -- .####...
                when x"31" & "0101" => d <= "00011000"; -- ...##...
                when x"31" & "0110" => d <= "00011000"; -- ...##...
                when x"31" & "0111" => d <= "00011000"; -- ...##...
                when x"31" & "1000" => d <= "00011000"; -- ...##...
                when x"31" & "1001" => d <= "00011000"; -- ...##...
                when x"31" & "1010" => d <= "00011000"; -- ...##...
                when x"31" & "1011" => d <= "01111110"; -- .######.
                when x"31" & "1100" => d <= "00000000"; -- ........
                when x"31" & "1101" => d <= "00000000"; -- ........
                when x"31" & "1110" => d <= "00000000"; -- ........
                when x"31" & "1111" => d <= "00000000"; -- ........

                when x"32" & "0000" => d <= "00000000"; -- ........
                when x"32" & "0001" => d <= "00000000"; -- ........
                when x"32" & "0010" => d <= "01111100"; -- .#####..
                when x"32" & "0011" => d <= "11000110"; -- ##...##.
                when x"32" & "0100" => d <= "00000110"; -- .....##.
                when x"32" & "0101" => d <= "00001100"; -- ....##..
                when x"32" & "0110" => d <= "00011000"; -- ...##...
                when x"32" & "0111" => d <= "00110000"; -- ..##....
                when x"32" & "1000" => d <= "01100000"; -- .##.....
                when x"32" & "1001" => d <= "11000000"; -- ##......
                when x"32" & "1010" => d <= "11000110"; -- ##...##.
                when x"32" & "1011" => d <= "11111110"; -- #######.
                when x"32" & "1100" => d <= "00000000"; -- ........
                when x"32" & "1101" => d <= "00000000"; -- ........
                when x"32" & "1110" => d <= "00000000"; -- ........
                when x"32" & "1111" => d <= "00000000"; -- ........

                when x"33" & "0000" => d <= "00000000"; -- ........
                when x"33" & "0001" => d <= "00000000"; -- ........
                when x"33" & "0010" => d <= "01111100"; -- .#####..
                when x"33" & "0011" => d <= "11000110"; -- ##...##.
                when x"33" & "0100" => d <= "00000110"; -- .....##.
                when x"33" & "0101" => d <= "00000110"; -- .....##.
                when x"33" & "0110" => d <= "00111100"; -- ..####..
                when x"33" & "0111" => d <= "00000110"; -- .....##.
                when x"33" & "1000" => d <= "00000110"; -- .....##.
                when x"33" & "1001" => d <= "00000110"; -- .....##.
                when x"33" & "1010" => d <= "11000110"; -- ##...##.
                when x"33" & "1011" => d <= "01111100"; -- .#####..
                when x"33" & "1100" => d <= "00000000"; -- ........
                when x"33" & "1101" => d <= "00000000"; -- ........
                when x"33" & "1110" => d <= "00000000"; -- ........
                when x"33" & "1111" => d <= "00000000"; -- ........

                when x"34" & "0000" => d <= "00000000"; -- ........
                when x"34" & "0001" => d <= "00000000"; -- ........
                when x"34" & "0010" => d <= "00001100"; -- ....##..
                when x"34" & "0011" => d <= "00011100"; -- ...###..
                when x"34" & "0100" => d <= "00111100"; -- ..####..
                when x"34" & "0101" => d <= "01101100"; -- .##.##..
                when x"34" & "0110" => d <= "11001100"; -- ##..##..
                when x"34" & "0111" => d <= "11111110"; -- #######.
                when x"34" & "1000" => d <= "00001100"; -- ....##..
                when x"34" & "1001" => d <= "00001100"; -- ....##..
                when x"34" & "1010" => d <= "00001100"; -- ....##..
                when x"34" & "1011" => d <= "00011110"; -- ...####.
                when x"34" & "1100" => d <= "00000000"; -- ........
                when x"34" & "1101" => d <= "00000000"; -- ........
                when x"34" & "1110" => d <= "00000000"; -- ........
                when x"34" & "1111" => d <= "00000000"; -- ........

                when x"35" & "0000" => d <= "00000000"; -- ........
                when x"35" & "0001" => d <= "00000000"; -- ........
                when x"35" & "0010" => d <= "11111110"; -- #######.
                when x"35" & "0011" => d <= "11000000"; -- ##......
                when x"35" & "0100" => d <= "11000000"; -- ##......
                when x"35" & "0101" => d <= "11000000"; -- ##......
                when x"35" & "0110" => d <= "11111100"; -- ######..
                when x"35" & "0111" => d <= "00000110"; -- .....##.
                when x"35" & "1000" => d <= "00000110"; -- .....##.
                when x"35" & "1001" => d <= "00000110"; -- .....##.
                when x"35" & "1010" => d <= "11000110"; -- ##...##.
                when x"35" & "1011" => d <= "01111100"; -- .#####..
                when x"35" & "1100" => d <= "00000000"; -- ........
                when x"35" & "1101" => d <= "00000000"; -- ........
                when x"35" & "1110" => d <= "00000000"; -- ........
                when x"35" & "1111" => d <= "00000000"; -- ........

                when x"36" & "0000" => d <= "00000000"; -- ........
                when x"36" & "0001" => d <= "00000000"; -- ........
                when x"36" & "0010" => d <= "00111000"; -- ..###...
                when x"36" & "0011" => d <= "01100000"; -- .##.....
                when x"36" & "0100" => d <= "11000000"; -- ##......
                when x"36" & "0101" => d <= "11000000"; -- ##......
                when x"36" & "0110" => d <= "11111100"; -- ######..
                when x"36" & "0111" => d <= "11000110"; -- ##...##.
                when x"36" & "1000" => d <= "11000110"; -- ##...##.
                when x"36" & "1001" => d <= "11000110"; -- ##...##.
                when x"36" & "1010" => d <= "11000110"; -- ##...##.
                when x"36" & "1011" => d <= "01111100"; -- .#####..
                when x"36" & "1100" => d <= "00000000"; -- ........
                when x"36" & "1101" => d <= "00000000"; -- ........
                when x"36" & "1110" => d <= "00000000"; -- ........
                when x"36" & "1111" => d <= "00000000"; -- ........

                when x"37" & "0000" => d <= "00000000"; -- ........
                when x"37" & "0001" => d <= "00000000"; -- ........
                when x"37" & "0010" => d <= "11111110"; -- #######.
                when x"37" & "0011" => d <= "11000110"; -- ##...##.
                when x"37" & "0100" => d <= "00000110"; -- .....##.
                when x"37" & "0101" => d <= "00000110"; -- .....##.
                when x"37" & "0110" => d <= "00001100"; -- ....##..
                when x"37" & "0111" => d <= "00011000"; -- ...##...
                when x"37" & "1000" => d <= "00110000"; -- ..##....
                when x"37" & "1001" => d <= "00110000"; -- ..##....
                when x"37" & "1010" => d <= "00110000"; -- ..##....
                when x"37" & "1011" => d <= "00110000"; -- ..##....
                when x"37" & "1100" => d <= "00000000"; -- ........
                when x"37" & "1101" => d <= "00000000"; -- ........
                when x"37" & "1110" => d <= "00000000"; -- ........
                when x"37" & "1111" => d <= "00000000"; -- ........

                when x"38" & "0000" => d <= "00000000"; -- ........
                when x"38" & "0001" => d <= "00000000"; -- ........
                when x"38" & "0010" => d <= "01111100"; -- .#####..
                when x"38" & "0011" => d <= "11000110"; -- ##...##.
                when x"38" & "0100" => d <= "11000110"; -- ##...##.
                when x"38" & "0101" => d <= "11000110"; -- ##...##.
                when x"38" & "0110" => d <= "01111100"; -- .#####..
                when x"38" & "0111" => d <= "11000110"; -- ##...##.
                when x"38" & "1000" => d <= "11000110"; -- ##...##.
                when x"38" & "1001" => d <= "11000110"; -- ##...##.
                when x"38" & "1010" => d <= "11000110"; -- ##...##.
                when x"38" & "1011" => d <= "01111100"; -- .#####..
                when x"38" & "1100" => d <= "00000000"; -- ........
                when x"38" & "1101" => d <= "00000000"; -- ........
                when x"38" & "1110" => d <= "00000000"; -- ........
                when x"38" & "1111" => d <= "00000000"; -- ........

                when x"39" & "0000" => d <= "00000000"; -- ........
                when x"39" & "0001" => d <= "00000000"; -- ........
                when x"39" & "0010" => d <= "01111100"; -- .#####..
                when x"39" & "0011" => d <= "11000110"; -- ##...##.
                when x"39" & "0100" => d <= "11000110"; -- ##...##.
                when x"39" & "0101" => d <= "11000110"; -- ##...##.
                when x"39" & "0110" => d <= "01111110"; -- .######.
                when x"39" & "0111" => d <= "00000110"; -- .....##.
                when x"39" & "1000" => d <= "00000110"; -- .....##.
                when x"39" & "1001" => d <= "00000110"; -- .....##.
                when x"39" & "1010" => d <= "00001100"; -- ....##..
                when x"39" & "1011" => d <= "01111000"; -- .####...
                when x"39" & "1100" => d <= "00000000"; -- ........
                when x"39" & "1101" => d <= "00000000"; -- ........
                when x"39" & "1110" => d <= "00000000"; -- ........
                when x"39" & "1111" => d <= "00000000"; -- ........

                when x"3a" & "0000" => d <= "00000000"; -- ........
                when x"3a" & "0001" => d <= "00000000"; -- ........
                when x"3a" & "0010" => d <= "00000000"; -- ........
                when x"3a" & "0011" => d <= "00000000"; -- ........
                when x"3a" & "0100" => d <= "00011000"; -- ...##...
                when x"3a" & "0101" => d <= "00011000"; -- ...##...
                when x"3a" & "0110" => d <= "00000000"; -- ........
                when x"3a" & "0111" => d <= "00000000"; -- ........
                when x"3a" & "1000" => d <= "00000000"; -- ........
                when x"3a" & "1001" => d <= "00011000"; -- ...##...
                when x"3a" & "1010" => d <= "00011000"; -- ...##...
                when x"3a" & "1011" => d <= "00000000"; -- ........
                when x"3a" & "1100" => d <= "00000000"; -- ........
                when x"3a" & "1101" => d <= "00000000"; -- ........
                when x"3a" & "1110" => d <= "00000000"; -- ........
                when x"3a" & "1111" => d <= "00000000"; -- ........

                when x"3b" & "0000" => d <= "00000000"; -- ........
                when x"3b" & "0001" => d <= "00000000"; -- ........
                when x"3b" & "0010" => d <= "00000000"; -- ........
                when x"3b" & "0011" => d <= "00000000"; -- ........
                when x"3b" & "0100" => d <= "00011000"; -- ...##...
                when x"3b" & "0101" => d <= "00011000"; -- ...##...
                when x"3b" & "0110" => d <= "00000000"; -- ........
                when x"3b" & "0111" => d <= "00000000"; -- ........
                when x"3b" & "1000" => d <= "00000000"; -- ........
                when x"3b" & "1001" => d <= "00011000"; -- ...##...
                when x"3b" & "1010" => d <= "00011000"; -- ...##...
                when x"3b" & "1011" => d <= "00110000"; -- ..##....
                when x"3b" & "1100" => d <= "00000000"; -- ........
                when x"3b" & "1101" => d <= "00000000"; -- ........
                when x"3b" & "1110" => d <= "00000000"; -- ........
                when x"3b" & "1111" => d <= "00000000"; -- ........

                when x"3c" & "0000" => d <= "00000000"; -- ........
                when x"3c" & "0001" => d <= "00000000"; -- ........
                when x"3c" & "0010" => d <= "00000000"; -- ........
                when x"3c" & "0011" => d <= "00000110"; -- .....##.
                when x"3c" & "0100" => d <= "00001100"; -- ....##..
                when x"3c" & "0101" => d <= "00011000"; -- ...##...
                when x"3c" & "0110" => d <= "00110000"; -- ..##....
                when x"3c" & "0111" => d <= "01100000"; -- .##.....
                when x"3c" & "1000" => d <= "00110000"; -- ..##....
                when x"3c" & "1001" => d <= "00011000"; -- ...##...
                when x"3c" & "1010" => d <= "00001100"; -- ....##..
                when x"3c" & "1011" => d <= "00000110"; -- .....##.
                when x"3c" & "1100" => d <= "00000000"; -- ........
                when x"3c" & "1101" => d <= "00000000"; -- ........
                when x"3c" & "1110" => d <= "00000000"; -- ........
                when x"3c" & "1111" => d <= "00000000"; -- ........

                when x"3d" & "0000" => d <= "00000000"; -- ........
                when x"3d" & "0001" => d <= "00000000"; -- ........
                when x"3d" & "0010" => d <= "00000000"; -- ........
                when x"3d" & "0011" => d <= "00000000"; -- ........
                when x"3d" & "0100" => d <= "00000000"; -- ........
                when x"3d" & "0101" => d <= "01111110"; -- .######.
                when x"3d" & "0110" => d <= "00000000"; -- ........
                when x"3d" & "0111" => d <= "00000000"; -- ........
                when x"3d" & "1000" => d <= "01111110"; -- .######.
                when x"3d" & "1001" => d <= "00000000"; -- ........
                when x"3d" & "1010" => d <= "00000000"; -- ........
                when x"3d" & "1011" => d <= "00000000"; -- ........
                when x"3d" & "1100" => d <= "00000000"; -- ........
                when x"3d" & "1101" => d <= "00000000"; -- ........
                when x"3d" & "1110" => d <= "00000000"; -- ........
                when x"3d" & "1111" => d <= "00000000"; -- ........

                when x"3e" & "0000" => d <= "00000000"; -- ........
                when x"3e" & "0001" => d <= "00000000"; -- ........
                when x"3e" & "0010" => d <= "00000000"; -- ........
                when x"3e" & "0011" => d <= "01100000"; -- .##.....
                when x"3e" & "0100" => d <= "00110000"; -- ..##....
                when x"3e" & "0101" => d <= "00011000"; -- ...##...
                when x"3e" & "0110" => d <= "00001100"; -- ....##..
                when x"3e" & "0111" => d <= "00000110"; -- .....##.
                when x"3e" & "1000" => d <= "00001100"; -- ....##..
                when x"3e" & "1001" => d <= "00011000"; -- ...##...
                when x"3e" & "1010" => d <= "00110000"; -- ..##....
                when x"3e" & "1011" => d <= "01100000"; -- .##.....
                when x"3e" & "1100" => d <= "00000000"; -- ........
                when x"3e" & "1101" => d <= "00000000"; -- ........
                when x"3e" & "1110" => d <= "00000000"; -- ........
                when x"3e" & "1111" => d <= "00000000"; -- ........

                when x"3f" & "0000" => d <= "00000000"; -- ........
                when x"3f" & "0001" => d <= "00000000"; -- ........
                when x"3f" & "0010" => d <= "01111100"; -- .#####..
                when x"3f" & "0011" => d <= "11000110"; -- ##...##.
                when x"3f" & "0100" => d <= "11000110"; -- ##...##.
                when x"3f" & "0101" => d <= "00001100"; -- ....##..
                when x"3f" & "0110" => d <= "00011000"; -- ...##...
                when x"3f" & "0111" => d <= "00011000"; -- ...##...
                when x"3f" & "1000" => d <= "00011000"; -- ...##...
                when x"3f" & "1001" => d <= "00000000"; -- ........
                when x"3f" & "1010" => d <= "00011000"; -- ...##...
                when x"3f" & "1011" => d <= "00011000"; -- ...##...
                when x"3f" & "1100" => d <= "00000000"; -- ........
                when x"3f" & "1101" => d <= "00000000"; -- ........
                when x"3f" & "1110" => d <= "00000000"; -- ........
                when x"3f" & "1111" => d <= "00000000"; -- ........

                when x"40" & "0000" => d <= "00000000"; -- ........
                when x"40" & "0001" => d <= "00000000"; -- ........
                when x"40" & "0010" => d <= "00000000"; -- ........
                when x"40" & "0011" => d <= "01111100"; -- .#####..
                when x"40" & "0100" => d <= "11000110"; -- ##...##.
                when x"40" & "0101" => d <= "11000110"; -- ##...##.
                when x"40" & "0110" => d <= "11011110"; -- ##.####.
                when x"40" & "0111" => d <= "11011110"; -- ##.####.
                when x"40" & "1000" => d <= "11011110"; -- ##.####.
                when x"40" & "1001" => d <= "11011100"; -- ##.###..
                when x"40" & "1010" => d <= "11000000"; -- ##......
                when x"40" & "1011" => d <= "01111100"; -- .#####..
                when x"40" & "1100" => d <= "00000000"; -- ........
                when x"40" & "1101" => d <= "00000000"; -- ........
                when x"40" & "1110" => d <= "00000000"; -- ........
                when x"40" & "1111" => d <= "00000000"; -- ........

                when x"41" & "0000" => d <= "00000000"; -- ........
                when x"41" & "0001" => d <= "00000000"; -- ........
                when x"41" & "0010" => d <= "00010000"; -- ...#....
                when x"41" & "0011" => d <= "00111000"; -- ..###...
                when x"41" & "0100" => d <= "01101100"; -- .##.##..
                when x"41" & "0101" => d <= "11000110"; -- ##...##.
                when x"41" & "0110" => d <= "11000110"; -- ##...##.
                when x"41" & "0111" => d <= "11111110"; -- #######.
                when x"41" & "1000" => d <= "11000110"; -- ##...##.
                when x"41" & "1001" => d <= "11000110"; -- ##...##.
                when x"41" & "1010" => d <= "11000110"; -- ##...##.
                when x"41" & "1011" => d <= "11000110"; -- ##...##.
                when x"41" & "1100" => d <= "00000000"; -- ........
                when x"41" & "1101" => d <= "00000000"; -- ........
                when x"41" & "1110" => d <= "00000000"; -- ........
                when x"41" & "1111" => d <= "00000000"; -- ........

                when x"42" & "0000" => d <= "00000000"; -- ........
                when x"42" & "0001" => d <= "00000000"; -- ........
                when x"42" & "0010" => d <= "11111100"; -- ######..
                when x"42" & "0011" => d <= "01100110"; -- .##..##.
                when x"42" & "0100" => d <= "01100110"; -- .##..##.
                when x"42" & "0101" => d <= "01100110"; -- .##..##.
                when x"42" & "0110" => d <= "01111100"; -- .#####..
                when x"42" & "0111" => d <= "01100110"; -- .##..##.
                when x"42" & "1000" => d <= "01100110"; -- .##..##.
                when x"42" & "1001" => d <= "01100110"; -- .##..##.
                when x"42" & "1010" => d <= "01100110"; -- .##..##.
                when x"42" & "1011" => d <= "11111100"; -- ######..
                when x"42" & "1100" => d <= "00000000"; -- ........
                when x"42" & "1101" => d <= "00000000"; -- ........
                when x"42" & "1110" => d <= "00000000"; -- ........
                when x"42" & "1111" => d <= "00000000"; -- ........

                when x"43" & "0000" => d <= "00000000"; -- ........
                when x"43" & "0001" => d <= "00000000"; -- ........
                when x"43" & "0010" => d <= "00111100"; -- ..####..
                when x"43" & "0011" => d <= "01100110"; -- .##..##.
                when x"43" & "0100" => d <= "11000010"; -- ##....#.
                when x"43" & "0101" => d <= "11000000"; -- ##......
                when x"43" & "0110" => d <= "11000000"; -- ##......
                when x"43" & "0111" => d <= "11000000"; -- ##......
                when x"43" & "1000" => d <= "11000000"; -- ##......
                when x"43" & "1001" => d <= "11000010"; -- ##....#.
                when x"43" & "1010" => d <= "01100110"; -- .##..##.
                when x"43" & "1011" => d <= "00111100"; -- ..####..
                when x"43" & "1100" => d <= "00000000"; -- ........
                when x"43" & "1101" => d <= "00000000"; -- ........
                when x"43" & "1110" => d <= "00000000"; -- ........
                when x"43" & "1111" => d <= "00000000"; -- ........

                when x"44" & "0000" => d <= "00000000"; -- ........
                when x"44" & "0001" => d <= "00000000"; -- ........
                when x"44" & "0010" => d <= "11111000"; -- #####...
                when x"44" & "0011" => d <= "01101100"; -- .##.##..
                when x"44" & "0100" => d <= "01100110"; -- .##..##.
                when x"44" & "0101" => d <= "01100110"; -- .##..##.
                when x"44" & "0110" => d <= "01100110"; -- .##..##.
                when x"44" & "0111" => d <= "01100110"; -- .##..##.
                when x"44" & "1000" => d <= "01100110"; -- .##..##.
                when x"44" & "1001" => d <= "01100110"; -- .##..##.
                when x"44" & "1010" => d <= "01101100"; -- .##.##..
                when x"44" & "1011" => d <= "11111000"; -- #####...
                when x"44" & "1100" => d <= "00000000"; -- ........
                when x"44" & "1101" => d <= "00000000"; -- ........
                when x"44" & "1110" => d <= "00000000"; -- ........
                when x"44" & "1111" => d <= "00000000"; -- ........

                when x"45" & "0000" => d <= "00000000"; -- ........
                when x"45" & "0001" => d <= "00000000"; -- ........
                when x"45" & "0010" => d <= "11111110"; -- #######.
                when x"45" & "0011" => d <= "01100110"; -- .##..##.
                when x"45" & "0100" => d <= "01100010"; -- .##...#.
                when x"45" & "0101" => d <= "01101000"; -- .##.#...
                when x"45" & "0110" => d <= "01111000"; -- .####...
                when x"45" & "0111" => d <= "01101000"; -- .##.#...
                when x"45" & "1000" => d <= "01100000"; -- .##.....
                when x"45" & "1001" => d <= "01100010"; -- .##...#.
                when x"45" & "1010" => d <= "01100110"; -- .##..##.
                when x"45" & "1011" => d <= "11111110"; -- #######.
                when x"45" & "1100" => d <= "00000000"; -- ........
                when x"45" & "1101" => d <= "00000000"; -- ........
                when x"45" & "1110" => d <= "00000000"; -- ........
                when x"45" & "1111" => d <= "00000000"; -- ........

                when x"46" & "0000" => d <= "00000000"; -- ........
                when x"46" & "0001" => d <= "00000000"; -- ........
                when x"46" & "0010" => d <= "11111110"; -- #######.
                when x"46" & "0011" => d <= "01100110"; -- .##..##.
                when x"46" & "0100" => d <= "01100010"; -- .##...#.
                when x"46" & "0101" => d <= "01101000"; -- .##.#...
                when x"46" & "0110" => d <= "01111000"; -- .####...
                when x"46" & "0111" => d <= "01101000"; -- .##.#...
                when x"46" & "1000" => d <= "01100000"; -- .##.....
                when x"46" & "1001" => d <= "01100000"; -- .##.....
                when x"46" & "1010" => d <= "01100000"; -- .##.....
                when x"46" & "1011" => d <= "11110000"; -- ####....
                when x"46" & "1100" => d <= "00000000"; -- ........
                when x"46" & "1101" => d <= "00000000"; -- ........
                when x"46" & "1110" => d <= "00000000"; -- ........
                when x"46" & "1111" => d <= "00000000"; -- ........

                when x"47" & "0000" => d <= "00000000"; -- ........
                when x"47" & "0001" => d <= "00000000"; -- ........
                when x"47" & "0010" => d <= "00111100"; -- ..####..
                when x"47" & "0011" => d <= "01100110"; -- .##..##.
                when x"47" & "0100" => d <= "11000010"; -- ##....#.
                when x"47" & "0101" => d <= "11000000"; -- ##......
                when x"47" & "0110" => d <= "11000000"; -- ##......
                when x"47" & "0111" => d <= "11011110"; -- ##.####.
                when x"47" & "1000" => d <= "11000110"; -- ##...##.
                when x"47" & "1001" => d <= "11000110"; -- ##...##.
                when x"47" & "1010" => d <= "01100110"; -- .##..##.
                when x"47" & "1011" => d <= "00111010"; -- ..###.#.
                when x"47" & "1100" => d <= "00000000"; -- ........
                when x"47" & "1101" => d <= "00000000"; -- ........
                when x"47" & "1110" => d <= "00000000"; -- ........
                when x"47" & "1111" => d <= "00000000"; -- ........

                when x"48" & "0000" => d <= "00000000"; -- ........
                when x"48" & "0001" => d <= "00000000"; -- ........
                when x"48" & "0010" => d <= "11000110"; -- ##...##.
                when x"48" & "0011" => d <= "11000110"; -- ##...##.
                when x"48" & "0100" => d <= "11000110"; -- ##...##.
                when x"48" & "0101" => d <= "11000110"; -- ##...##.
                when x"48" & "0110" => d <= "11111110"; -- #######.
                when x"48" & "0111" => d <= "11000110"; -- ##...##.
                when x"48" & "1000" => d <= "11000110"; -- ##...##.
                when x"48" & "1001" => d <= "11000110"; -- ##...##.
                when x"48" & "1010" => d <= "11000110"; -- ##...##.
                when x"48" & "1011" => d <= "11000110"; -- ##...##.
                when x"48" & "1100" => d <= "00000000"; -- ........
                when x"48" & "1101" => d <= "00000000"; -- ........
                when x"48" & "1110" => d <= "00000000"; -- ........
                when x"48" & "1111" => d <= "00000000"; -- ........

                when x"49" & "0000" => d <= "00000000"; -- ........
                when x"49" & "0001" => d <= "00000000"; -- ........
                when x"49" & "0010" => d <= "00111100"; -- ..####..
                when x"49" & "0011" => d <= "00011000"; -- ...##...
                when x"49" & "0100" => d <= "00011000"; -- ...##...
                when x"49" & "0101" => d <= "00011000"; -- ...##...
                when x"49" & "0110" => d <= "00011000"; -- ...##...
                when x"49" & "0111" => d <= "00011000"; -- ...##...
                when x"49" & "1000" => d <= "00011000"; -- ...##...
                when x"49" & "1001" => d <= "00011000"; -- ...##...
                when x"49" & "1010" => d <= "00011000"; -- ...##...
                when x"49" & "1011" => d <= "00111100"; -- ..####..
                when x"49" & "1100" => d <= "00000000"; -- ........
                when x"49" & "1101" => d <= "00000000"; -- ........
                when x"49" & "1110" => d <= "00000000"; -- ........
                when x"49" & "1111" => d <= "00000000"; -- ........

                when x"4a" & "0000" => d <= "00000000"; -- ........
                when x"4a" & "0001" => d <= "00000000"; -- ........
                when x"4a" & "0010" => d <= "00011110"; -- ...####.
                when x"4a" & "0011" => d <= "00001100"; -- ....##..
                when x"4a" & "0100" => d <= "00001100"; -- ....##..
                when x"4a" & "0101" => d <= "00001100"; -- ....##..
                when x"4a" & "0110" => d <= "00001100"; -- ....##..
                when x"4a" & "0111" => d <= "00001100"; -- ....##..
                when x"4a" & "1000" => d <= "11001100"; -- ##..##..
                when x"4a" & "1001" => d <= "11001100"; -- ##..##..
                when x"4a" & "1010" => d <= "11001100"; -- ##..##..
                when x"4a" & "1011" => d <= "01111000"; -- .####...
                when x"4a" & "1100" => d <= "00000000"; -- ........
                when x"4a" & "1101" => d <= "00000000"; -- ........
                when x"4a" & "1110" => d <= "00000000"; -- ........
                when x"4a" & "1111" => d <= "00000000"; -- ........

                when x"4b" & "0000" => d <= "00000000"; -- ........
                when x"4b" & "0001" => d <= "00000000"; -- ........
                when x"4b" & "0010" => d <= "11100110"; -- ###..##.
                when x"4b" & "0011" => d <= "01100110"; -- .##..##.
                when x"4b" & "0100" => d <= "01100110"; -- .##..##.
                when x"4b" & "0101" => d <= "01101100"; -- .##.##..
                when x"4b" & "0110" => d <= "01111000"; -- .####...
                when x"4b" & "0111" => d <= "01111000"; -- .####...
                when x"4b" & "1000" => d <= "01101100"; -- .##.##..
                when x"4b" & "1001" => d <= "01100110"; -- .##..##.
                when x"4b" & "1010" => d <= "01100110"; -- .##..##.
                when x"4b" & "1011" => d <= "11100110"; -- ###..##.
                when x"4b" & "1100" => d <= "00000000"; -- ........
                when x"4b" & "1101" => d <= "00000000"; -- ........
                when x"4b" & "1110" => d <= "00000000"; -- ........
                when x"4b" & "1111" => d <= "00000000"; -- ........

                when x"4c" & "0000" => d <= "00000000"; -- ........
                when x"4c" & "0001" => d <= "00000000"; -- ........
                when x"4c" & "0010" => d <= "11110000"; -- ####....
                when x"4c" & "0011" => d <= "01100000"; -- .##.....
                when x"4c" & "0100" => d <= "01100000"; -- .##.....
                when x"4c" & "0101" => d <= "01100000"; -- .##.....
                when x"4c" & "0110" => d <= "01100000"; -- .##.....
                when x"4c" & "0111" => d <= "01100000"; -- .##.....
                when x"4c" & "1000" => d <= "01100000"; -- .##.....
                when x"4c" & "1001" => d <= "01100010"; -- .##...#.
                when x"4c" & "1010" => d <= "01100110"; -- .##..##.
                when x"4c" & "1011" => d <= "11111110"; -- #######.
                when x"4c" & "1100" => d <= "00000000"; -- ........
                when x"4c" & "1101" => d <= "00000000"; -- ........
                when x"4c" & "1110" => d <= "00000000"; -- ........
                when x"4c" & "1111" => d <= "00000000"; -- ........

                when x"4d" & "0000" => d <= "00000000"; -- ........
                when x"4d" & "0001" => d <= "00000000"; -- ........
                when x"4d" & "0010" => d <= "11000110"; -- ##...##.
                when x"4d" & "0011" => d <= "11101110"; -- ###.###.
                when x"4d" & "0100" => d <= "11111110"; -- #######.
                when x"4d" & "0101" => d <= "11111110"; -- #######.
                when x"4d" & "0110" => d <= "11010110"; -- ##.#.##.
                when x"4d" & "0111" => d <= "11000110"; -- ##...##.
                when x"4d" & "1000" => d <= "11000110"; -- ##...##.
                when x"4d" & "1001" => d <= "11000110"; -- ##...##.
                when x"4d" & "1010" => d <= "11000110"; -- ##...##.
                when x"4d" & "1011" => d <= "11000110"; -- ##...##.
                when x"4d" & "1100" => d <= "00000000"; -- ........
                when x"4d" & "1101" => d <= "00000000"; -- ........
                when x"4d" & "1110" => d <= "00000000"; -- ........
                when x"4d" & "1111" => d <= "00000000"; -- ........

                when x"4e" & "0000" => d <= "00000000"; -- ........
                when x"4e" & "0001" => d <= "00000000"; -- ........
                when x"4e" & "0010" => d <= "11000110"; -- ##...##.
                when x"4e" & "0011" => d <= "11100110"; -- ###..##.
                when x"4e" & "0100" => d <= "11110110"; -- ####.##.
                when x"4e" & "0101" => d <= "11111110"; -- #######.
                when x"4e" & "0110" => d <= "11011110"; -- ##.####.
                when x"4e" & "0111" => d <= "11001110"; -- ##..###.
                when x"4e" & "1000" => d <= "11000110"; -- ##...##.
                when x"4e" & "1001" => d <= "11000110"; -- ##...##.
                when x"4e" & "1010" => d <= "11000110"; -- ##...##.
                when x"4e" & "1011" => d <= "11000110"; -- ##...##.
                when x"4e" & "1100" => d <= "00000000"; -- ........
                when x"4e" & "1101" => d <= "00000000"; -- ........
                when x"4e" & "1110" => d <= "00000000"; -- ........
                when x"4e" & "1111" => d <= "00000000"; -- ........

                when x"4f" & "0000" => d <= "00000000"; -- ........
                when x"4f" & "0001" => d <= "00000000"; -- ........
                when x"4f" & "0010" => d <= "01111100"; -- .#####..
                when x"4f" & "0011" => d <= "11000110"; -- ##...##.
                when x"4f" & "0100" => d <= "11000110"; -- ##...##.
                when x"4f" & "0101" => d <= "11000110"; -- ##...##.
                when x"4f" & "0110" => d <= "11000110"; -- ##...##.
                when x"4f" & "0111" => d <= "11000110"; -- ##...##.
                when x"4f" & "1000" => d <= "11000110"; -- ##...##.
                when x"4f" & "1001" => d <= "11000110"; -- ##...##.
                when x"4f" & "1010" => d <= "11000110"; -- ##...##.
                when x"4f" & "1011" => d <= "01111100"; -- .#####..
                when x"4f" & "1100" => d <= "00000000"; -- ........
                when x"4f" & "1101" => d <= "00000000"; -- ........
                when x"4f" & "1110" => d <= "00000000"; -- ........
                when x"4f" & "1111" => d <= "00000000"; -- ........

                when x"50" & "0000" => d <= "00000000"; -- ........
                when x"50" & "0001" => d <= "00000000"; -- ........
                when x"50" & "0010" => d <= "11111100"; -- ######..
                when x"50" & "0011" => d <= "01100110"; -- .##..##.
                when x"50" & "0100" => d <= "01100110"; -- .##..##.
                when x"50" & "0101" => d <= "01100110"; -- .##..##.
                when x"50" & "0110" => d <= "01111100"; -- .#####..
                when x"50" & "0111" => d <= "01100000"; -- .##.....
                when x"50" & "1000" => d <= "01100000"; -- .##.....
                when x"50" & "1001" => d <= "01100000"; -- .##.....
                when x"50" & "1010" => d <= "01100000"; -- .##.....
                when x"50" & "1011" => d <= "11110000"; -- ####....
                when x"50" & "1100" => d <= "00000000"; -- ........
                when x"50" & "1101" => d <= "00000000"; -- ........
                when x"50" & "1110" => d <= "00000000"; -- ........
                when x"50" & "1111" => d <= "00000000"; -- ........

                when x"51" & "0000" => d <= "00000000"; -- ........
                when x"51" & "0001" => d <= "00000000"; -- ........
                when x"51" & "0010" => d <= "01111100"; -- .#####..
                when x"51" & "0011" => d <= "11000110"; -- ##...##.
                when x"51" & "0100" => d <= "11000110"; -- ##...##.
                when x"51" & "0101" => d <= "11000110"; -- ##...##.
                when x"51" & "0110" => d <= "11000110"; -- ##...##.
                when x"51" & "0111" => d <= "11000110"; -- ##...##.
                when x"51" & "1000" => d <= "11000110"; -- ##...##.
                when x"51" & "1001" => d <= "11010110"; -- ##.#.##.
                when x"51" & "1010" => d <= "11011110"; -- ##.####.
                when x"51" & "1011" => d <= "01111100"; -- .#####..
                when x"51" & "1100" => d <= "00001100"; -- ....##..
                when x"51" & "1101" => d <= "00001110"; -- ....###.
                when x"51" & "1110" => d <= "00000000"; -- ........
                when x"51" & "1111" => d <= "00000000"; -- ........

                when x"52" & "0000" => d <= "00000000"; -- ........
                when x"52" & "0001" => d <= "00000000"; -- ........
                when x"52" & "0010" => d <= "11111100"; -- ######..
                when x"52" & "0011" => d <= "01100110"; -- .##..##.
                when x"52" & "0100" => d <= "01100110"; -- .##..##.
                when x"52" & "0101" => d <= "01100110"; -- .##..##.
                when x"52" & "0110" => d <= "01111100"; -- .#####..
                when x"52" & "0111" => d <= "01101100"; -- .##.##..
                when x"52" & "1000" => d <= "01100110"; -- .##..##.
                when x"52" & "1001" => d <= "01100110"; -- .##..##.
                when x"52" & "1010" => d <= "01100110"; -- .##..##.
                when x"52" & "1011" => d <= "11100110"; -- ###..##.
                when x"52" & "1100" => d <= "00000000"; -- ........
                when x"52" & "1101" => d <= "00000000"; -- ........
                when x"52" & "1110" => d <= "00000000"; -- ........
                when x"52" & "1111" => d <= "00000000"; -- ........

                when x"53" & "0000" => d <= "00000000"; -- ........
                when x"53" & "0001" => d <= "00000000"; -- ........
                when x"53" & "0010" => d <= "01111100"; -- .#####..
                when x"53" & "0011" => d <= "11000110"; -- ##...##.
                when x"53" & "0100" => d <= "11000110"; -- ##...##.
                when x"53" & "0101" => d <= "01100000"; -- .##.....
                when x"53" & "0110" => d <= "00111000"; -- ..###...
                when x"53" & "0111" => d <= "00001100"; -- ....##..
                when x"53" & "1000" => d <= "00000110"; -- .....##.
                when x"53" & "1001" => d <= "11000110"; -- ##...##.
                when x"53" & "1010" => d <= "11000110"; -- ##...##.
                when x"53" & "1011" => d <= "01111100"; -- .#####..
                when x"53" & "1100" => d <= "00000000"; -- ........
                when x"53" & "1101" => d <= "00000000"; -- ........
                when x"53" & "1110" => d <= "00000000"; -- ........
                when x"53" & "1111" => d <= "00000000"; -- ........

                when x"54" & "0000" => d <= "00000000"; -- ........
                when x"54" & "0001" => d <= "00000000"; -- ........
                when x"54" & "0010" => d <= "01111110"; -- .######.
                when x"54" & "0011" => d <= "01111110"; -- .######.
                when x"54" & "0100" => d <= "01011010"; -- .#.##.#.
                when x"54" & "0101" => d <= "00011000"; -- ...##...
                when x"54" & "0110" => d <= "00011000"; -- ...##...
                when x"54" & "0111" => d <= "00011000"; -- ...##...
                when x"54" & "1000" => d <= "00011000"; -- ...##...
                when x"54" & "1001" => d <= "00011000"; -- ...##...
                when x"54" & "1010" => d <= "00011000"; -- ...##...
                when x"54" & "1011" => d <= "00111100"; -- ..####..
                when x"54" & "1100" => d <= "00000000"; -- ........
                when x"54" & "1101" => d <= "00000000"; -- ........
                when x"54" & "1110" => d <= "00000000"; -- ........
                when x"54" & "1111" => d <= "00000000"; -- ........

                when x"55" & "0000" => d <= "00000000"; -- ........
                when x"55" & "0001" => d <= "00000000"; -- ........
                when x"55" & "0010" => d <= "11000110"; -- ##...##.
                when x"55" & "0011" => d <= "11000110"; -- ##...##.
                when x"55" & "0100" => d <= "11000110"; -- ##...##.
                when x"55" & "0101" => d <= "11000110"; -- ##...##.
                when x"55" & "0110" => d <= "11000110"; -- ##...##.
                when x"55" & "0111" => d <= "11000110"; -- ##...##.
                when x"55" & "1000" => d <= "11000110"; -- ##...##.
                when x"55" & "1001" => d <= "11000110"; -- ##...##.
                when x"55" & "1010" => d <= "11000110"; -- ##...##.
                when x"55" & "1011" => d <= "01111100"; -- .#####..
                when x"55" & "1100" => d <= "00000000"; -- ........
                when x"55" & "1101" => d <= "00000000"; -- ........
                when x"55" & "1110" => d <= "00000000"; -- ........
                when x"55" & "1111" => d <= "00000000"; -- ........

                when x"56" & "0000" => d <= "00000000"; -- ........
                when x"56" & "0001" => d <= "00000000"; -- ........
                when x"56" & "0010" => d <= "11000110"; -- ##...##.
                when x"56" & "0011" => d <= "11000110"; -- ##...##.
                when x"56" & "0100" => d <= "11000110"; -- ##...##.
                when x"56" & "0101" => d <= "11000110"; -- ##...##.
                when x"56" & "0110" => d <= "11000110"; -- ##...##.
                when x"56" & "0111" => d <= "11000110"; -- ##...##.
                when x"56" & "1000" => d <= "11000110"; -- ##...##.
                when x"56" & "1001" => d <= "01101100"; -- .##.##..
                when x"56" & "1010" => d <= "00111000"; -- ..###...
                when x"56" & "1011" => d <= "00010000"; -- ...#....
                when x"56" & "1100" => d <= "00000000"; -- ........
                when x"56" & "1101" => d <= "00000000"; -- ........
                when x"56" & "1110" => d <= "00000000"; -- ........
                when x"56" & "1111" => d <= "00000000"; -- ........

                when x"57" & "0000" => d <= "00000000"; -- ........
                when x"57" & "0001" => d <= "00000000"; -- ........
                when x"57" & "0010" => d <= "11000110"; -- ##...##.
                when x"57" & "0011" => d <= "11000110"; -- ##...##.
                when x"57" & "0100" => d <= "11000110"; -- ##...##.
                when x"57" & "0101" => d <= "11000110"; -- ##...##.
                when x"57" & "0110" => d <= "11010110"; -- ##.#.##.
                when x"57" & "0111" => d <= "11010110"; -- ##.#.##.
                when x"57" & "1000" => d <= "11010110"; -- ##.#.##.
                when x"57" & "1001" => d <= "11111110"; -- #######.
                when x"57" & "1010" => d <= "11101110"; -- ###.###.
                when x"57" & "1011" => d <= "01101100"; -- .##.##..
                when x"57" & "1100" => d <= "00000000"; -- ........
                when x"57" & "1101" => d <= "00000000"; -- ........
                when x"57" & "1110" => d <= "00000000"; -- ........
                when x"57" & "1111" => d <= "00000000"; -- ........

                when x"58" & "0000" => d <= "00000000"; -- ........
                when x"58" & "0001" => d <= "00000000"; -- ........
                when x"58" & "0010" => d <= "11000110"; -- ##...##.
                when x"58" & "0011" => d <= "11000110"; -- ##...##.
                when x"58" & "0100" => d <= "01101100"; -- .##.##..
                when x"58" & "0101" => d <= "01111100"; -- .#####..
                when x"58" & "0110" => d <= "00111000"; -- ..###...
                when x"58" & "0111" => d <= "00111000"; -- ..###...
                when x"58" & "1000" => d <= "01111100"; -- .#####..
                when x"58" & "1001" => d <= "01101100"; -- .##.##..
                when x"58" & "1010" => d <= "11000110"; -- ##...##.
                when x"58" & "1011" => d <= "11000110"; -- ##...##.
                when x"58" & "1100" => d <= "00000000"; -- ........
                when x"58" & "1101" => d <= "00000000"; -- ........
                when x"58" & "1110" => d <= "00000000"; -- ........
                when x"58" & "1111" => d <= "00000000"; -- ........

                when x"59" & "0000" => d <= "00000000"; -- ........
                when x"59" & "0001" => d <= "00000000"; -- ........
                when x"59" & "0010" => d <= "01100110"; -- .##..##.
                when x"59" & "0011" => d <= "01100110"; -- .##..##.
                when x"59" & "0100" => d <= "01100110"; -- .##..##.
                when x"59" & "0101" => d <= "01100110"; -- .##..##.
                when x"59" & "0110" => d <= "00111100"; -- ..####..
                when x"59" & "0111" => d <= "00011000"; -- ...##...
                when x"59" & "1000" => d <= "00011000"; -- ...##...
                when x"59" & "1001" => d <= "00011000"; -- ...##...
                when x"59" & "1010" => d <= "00011000"; -- ...##...
                when x"59" & "1011" => d <= "00111100"; -- ..####..
                when x"59" & "1100" => d <= "00000000"; -- ........
                when x"59" & "1101" => d <= "00000000"; -- ........
                when x"59" & "1110" => d <= "00000000"; -- ........
                when x"59" & "1111" => d <= "00000000"; -- ........

                when x"5a" & "0000" => d <= "00000000"; -- ........
                when x"5a" & "0001" => d <= "00000000"; -- ........
                when x"5a" & "0010" => d <= "11111110"; -- #######.
                when x"5a" & "0011" => d <= "11000110"; -- ##...##.
                when x"5a" & "0100" => d <= "10000110"; -- #....##.
                when x"5a" & "0101" => d <= "00001100"; -- ....##..
                when x"5a" & "0110" => d <= "00011000"; -- ...##...
                when x"5a" & "0111" => d <= "00110000"; -- ..##....
                when x"5a" & "1000" => d <= "01100000"; -- .##.....
                when x"5a" & "1001" => d <= "11000010"; -- ##....#.
                when x"5a" & "1010" => d <= "11000110"; -- ##...##.
                when x"5a" & "1011" => d <= "11111110"; -- #######.
                when x"5a" & "1100" => d <= "00000000"; -- ........
                when x"5a" & "1101" => d <= "00000000"; -- ........
                when x"5a" & "1110" => d <= "00000000"; -- ........
                when x"5a" & "1111" => d <= "00000000"; -- ........

                when x"5b" & "0000" => d <= "00000000"; -- ........
                when x"5b" & "0001" => d <= "00000000"; -- ........
                when x"5b" & "0010" => d <= "00111100"; -- ..####..
                when x"5b" & "0011" => d <= "00110000"; -- ..##....
                when x"5b" & "0100" => d <= "00110000"; -- ..##....
                when x"5b" & "0101" => d <= "00110000"; -- ..##....
                when x"5b" & "0110" => d <= "00110000"; -- ..##....
                when x"5b" & "0111" => d <= "00110000"; -- ..##....
                when x"5b" & "1000" => d <= "00110000"; -- ..##....
                when x"5b" & "1001" => d <= "00110000"; -- ..##....
                when x"5b" & "1010" => d <= "00110000"; -- ..##....
                when x"5b" & "1011" => d <= "00111100"; -- ..####..
                when x"5b" & "1100" => d <= "00000000"; -- ........
                when x"5b" & "1101" => d <= "00000000"; -- ........
                when x"5b" & "1110" => d <= "00000000"; -- ........
                when x"5b" & "1111" => d <= "00000000"; -- ........

                when x"5c" & "0000" => d <= "00000000"; -- ........
                when x"5c" & "0001" => d <= "00000000"; -- ........
                when x"5c" & "0010" => d <= "00000000"; -- ........
                when x"5c" & "0011" => d <= "10000000"; -- #.......
                when x"5c" & "0100" => d <= "11000000"; -- ##......
                when x"5c" & "0101" => d <= "11100000"; -- ###.....
                when x"5c" & "0110" => d <= "01110000"; -- .###....
                when x"5c" & "0111" => d <= "00111000"; -- ..###...
                when x"5c" & "1000" => d <= "00011100"; -- ...###..
                when x"5c" & "1001" => d <= "00001110"; -- ....###.
                when x"5c" & "1010" => d <= "00000110"; -- .....##.
                when x"5c" & "1011" => d <= "00000010"; -- ......#.
                when x"5c" & "1100" => d <= "00000000"; -- ........
                when x"5c" & "1101" => d <= "00000000"; -- ........
                when x"5c" & "1110" => d <= "00000000"; -- ........
                when x"5c" & "1111" => d <= "00000000"; -- ........

                when x"5d" & "0000" => d <= "00000000"; -- ........
                when x"5d" & "0001" => d <= "00000000"; -- ........
                when x"5d" & "0010" => d <= "00111100"; -- ..####..
                when x"5d" & "0011" => d <= "00001100"; -- ....##..
                when x"5d" & "0100" => d <= "00001100"; -- ....##..
                when x"5d" & "0101" => d <= "00001100"; -- ....##..
                when x"5d" & "0110" => d <= "00001100"; -- ....##..
                when x"5d" & "0111" => d <= "00001100"; -- ....##..
                when x"5d" & "1000" => d <= "00001100"; -- ....##..
                when x"5d" & "1001" => d <= "00001100"; -- ....##..
                when x"5d" & "1010" => d <= "00001100"; -- ....##..
                when x"5d" & "1011" => d <= "00111100"; -- ..####..
                when x"5d" & "1100" => d <= "00000000"; -- ........
                when x"5d" & "1101" => d <= "00000000"; -- ........
                when x"5d" & "1110" => d <= "00000000"; -- ........
                when x"5d" & "1111" => d <= "00000000"; -- ........

                when x"5e" & "0000" => d <= "00010000"; -- ...#....
                when x"5e" & "0001" => d <= "00111000"; -- ..###...
                when x"5e" & "0010" => d <= "01101100"; -- .##.##..
                when x"5e" & "0011" => d <= "11000110"; -- ##...##.
                when x"5e" & "0100" => d <= "00000000"; -- ........
                when x"5e" & "0101" => d <= "00000000"; -- ........
                when x"5e" & "0110" => d <= "00000000"; -- ........
                when x"5e" & "0111" => d <= "00000000"; -- ........
                when x"5e" & "1000" => d <= "00000000"; -- ........
                when x"5e" & "1001" => d <= "00000000"; -- ........
                when x"5e" & "1010" => d <= "00000000"; -- ........
                when x"5e" & "1011" => d <= "00000000"; -- ........
                when x"5e" & "1100" => d <= "00000000"; -- ........
                when x"5e" & "1101" => d <= "00000000"; -- ........
                when x"5e" & "1110" => d <= "00000000"; -- ........
                when x"5e" & "1111" => d <= "00000000"; -- ........

                when x"5f" & "0000" => d <= "00000000"; -- ........
                when x"5f" & "0001" => d <= "00000000"; -- ........
                when x"5f" & "0010" => d <= "00000000"; -- ........
                when x"5f" & "0011" => d <= "00000000"; -- ........
                when x"5f" & "0100" => d <= "00000000"; -- ........
                when x"5f" & "0101" => d <= "00000000"; -- ........
                when x"5f" & "0110" => d <= "00000000"; -- ........
                when x"5f" & "0111" => d <= "00000000"; -- ........
                when x"5f" & "1000" => d <= "00000000"; -- ........
                when x"5f" & "1001" => d <= "00000000"; -- ........
                when x"5f" & "1010" => d <= "00000000"; -- ........
                when x"5f" & "1011" => d <= "00000000"; -- ........
                when x"5f" & "1100" => d <= "00000000"; -- ........
                when x"5f" & "1101" => d <= "11111111"; -- ########
                when x"5f" & "1110" => d <= "00000000"; -- ........
                when x"5f" & "1111" => d <= "00000000"; -- ........

                when x"60" & "0000" => d <= "00110000"; -- ..##....
                when x"60" & "0001" => d <= "00110000"; -- ..##....
                when x"60" & "0010" => d <= "00011000"; -- ...##...
                when x"60" & "0011" => d <= "00000000"; -- ........
                when x"60" & "0100" => d <= "00000000"; -- ........
                when x"60" & "0101" => d <= "00000000"; -- ........
                when x"60" & "0110" => d <= "00000000"; -- ........
                when x"60" & "0111" => d <= "00000000"; -- ........
                when x"60" & "1000" => d <= "00000000"; -- ........
                when x"60" & "1001" => d <= "00000000"; -- ........
                when x"60" & "1010" => d <= "00000000"; -- ........
                when x"60" & "1011" => d <= "00000000"; -- ........
                when x"60" & "1100" => d <= "00000000"; -- ........
                when x"60" & "1101" => d <= "00000000"; -- ........
                when x"60" & "1110" => d <= "00000000"; -- ........
                when x"60" & "1111" => d <= "00000000"; -- ........

                when x"61" & "0000" => d <= "00000000"; -- ........
                when x"61" & "0001" => d <= "00000000"; -- ........
                when x"61" & "0010" => d <= "00000000"; -- ........
                when x"61" & "0011" => d <= "00000000"; -- ........
                when x"61" & "0100" => d <= "00000000"; -- ........
                when x"61" & "0101" => d <= "01111000"; -- .####...
                when x"61" & "0110" => d <= "00001100"; -- ....##..
                when x"61" & "0111" => d <= "01111100"; -- .#####..
                when x"61" & "1000" => d <= "11001100"; -- ##..##..
                when x"61" & "1001" => d <= "11001100"; -- ##..##..
                when x"61" & "1010" => d <= "11001100"; -- ##..##..
                when x"61" & "1011" => d <= "01110110"; -- .###.##.
                when x"61" & "1100" => d <= "00000000"; -- ........
                when x"61" & "1101" => d <= "00000000"; -- ........
                when x"61" & "1110" => d <= "00000000"; -- ........
                when x"61" & "1111" => d <= "00000000"; -- ........

                when x"62" & "0000" => d <= "00000000"; -- ........
                when x"62" & "0001" => d <= "00000000"; -- ........
                when x"62" & "0010" => d <= "11100000"; -- ###.....
                when x"62" & "0011" => d <= "01100000"; -- .##.....
                when x"62" & "0100" => d <= "01100000"; -- .##.....
                when x"62" & "0101" => d <= "01111000"; -- .####...
                when x"62" & "0110" => d <= "01101100"; -- .##.##..
                when x"62" & "0111" => d <= "01100110"; -- .##..##.
                when x"62" & "1000" => d <= "01100110"; -- .##..##.
                when x"62" & "1001" => d <= "01100110"; -- .##..##.
                when x"62" & "1010" => d <= "01100110"; -- .##..##.
                when x"62" & "1011" => d <= "01111100"; -- .#####..
                when x"62" & "1100" => d <= "00000000"; -- ........
                when x"62" & "1101" => d <= "00000000"; -- ........
                when x"62" & "1110" => d <= "00000000"; -- ........
                when x"62" & "1111" => d <= "00000000"; -- ........

                when x"63" & "0000" => d <= "00000000"; -- ........
                when x"63" & "0001" => d <= "00000000"; -- ........
                when x"63" & "0010" => d <= "00000000"; -- ........
                when x"63" & "0011" => d <= "00000000"; -- ........
                when x"63" & "0100" => d <= "00000000"; -- ........
                when x"63" & "0101" => d <= "01111100"; -- .#####..
                when x"63" & "0110" => d <= "11000110"; -- ##...##.
                when x"63" & "0111" => d <= "11000000"; -- ##......
                when x"63" & "1000" => d <= "11000000"; -- ##......
                when x"63" & "1001" => d <= "11000000"; -- ##......
                when x"63" & "1010" => d <= "11000110"; -- ##...##.
                when x"63" & "1011" => d <= "01111100"; -- .#####..
                when x"63" & "1100" => d <= "00000000"; -- ........
                when x"63" & "1101" => d <= "00000000"; -- ........
                when x"63" & "1110" => d <= "00000000"; -- ........
                when x"63" & "1111" => d <= "00000000"; -- ........

                when x"64" & "0000" => d <= "00000000"; -- ........
                when x"64" & "0001" => d <= "00000000"; -- ........
                when x"64" & "0010" => d <= "00011100"; -- ...###..
                when x"64" & "0011" => d <= "00001100"; -- ....##..
                when x"64" & "0100" => d <= "00001100"; -- ....##..
                when x"64" & "0101" => d <= "00111100"; -- ..####..
                when x"64" & "0110" => d <= "01101100"; -- .##.##..
                when x"64" & "0111" => d <= "11001100"; -- ##..##..
                when x"64" & "1000" => d <= "11001100"; -- ##..##..
                when x"64" & "1001" => d <= "11001100"; -- ##..##..
                when x"64" & "1010" => d <= "11001100"; -- ##..##..
                when x"64" & "1011" => d <= "01110110"; -- .###.##.
                when x"64" & "1100" => d <= "00000000"; -- ........
                when x"64" & "1101" => d <= "00000000"; -- ........
                when x"64" & "1110" => d <= "00000000"; -- ........
                when x"64" & "1111" => d <= "00000000"; -- ........

                when x"65" & "0000" => d <= "00000000"; -- ........
                when x"65" & "0001" => d <= "00000000"; -- ........
                when x"65" & "0010" => d <= "00000000"; -- ........
                when x"65" & "0011" => d <= "00000000"; -- ........
                when x"65" & "0100" => d <= "00000000"; -- ........
                when x"65" & "0101" => d <= "01111100"; -- .#####..
                when x"65" & "0110" => d <= "11000110"; -- ##...##.
                when x"65" & "0111" => d <= "11111110"; -- #######.
                when x"65" & "1000" => d <= "11000000"; -- ##......
                when x"65" & "1001" => d <= "11000000"; -- ##......
                when x"65" & "1010" => d <= "11000110"; -- ##...##.
                when x"65" & "1011" => d <= "01111100"; -- .#####..
                when x"65" & "1100" => d <= "00000000"; -- ........
                when x"65" & "1101" => d <= "00000000"; -- ........
                when x"65" & "1110" => d <= "00000000"; -- ........
                when x"65" & "1111" => d <= "00000000"; -- ........

                when x"66" & "0000" => d <= "00000000"; -- ........
                when x"66" & "0001" => d <= "00000000"; -- ........
                when x"66" & "0010" => d <= "00111000"; -- ..###...
                when x"66" & "0011" => d <= "01101100"; -- .##.##..
                when x"66" & "0100" => d <= "01100100"; -- .##..#..
                when x"66" & "0101" => d <= "01100000"; -- .##.....
                when x"66" & "0110" => d <= "11110000"; -- ####....
                when x"66" & "0111" => d <= "01100000"; -- .##.....
                when x"66" & "1000" => d <= "01100000"; -- .##.....
                when x"66" & "1001" => d <= "01100000"; -- .##.....
                when x"66" & "1010" => d <= "01100000"; -- .##.....
                when x"66" & "1011" => d <= "11110000"; -- ####....
                when x"66" & "1100" => d <= "00000000"; -- ........
                when x"66" & "1101" => d <= "00000000"; -- ........
                when x"66" & "1110" => d <= "00000000"; -- ........
                when x"66" & "1111" => d <= "00000000"; -- ........

                when x"67" & "0000" => d <= "00000000"; -- ........
                when x"67" & "0001" => d <= "00000000"; -- ........
                when x"67" & "0010" => d <= "00000000"; -- ........
                when x"67" & "0011" => d <= "00000000"; -- ........
                when x"67" & "0100" => d <= "00000000"; -- ........
                when x"67" & "0101" => d <= "01110110"; -- .###.##.
                when x"67" & "0110" => d <= "11001100"; -- ##..##..
                when x"67" & "0111" => d <= "11001100"; -- ##..##..
                when x"67" & "1000" => d <= "11001100"; -- ##..##..
                when x"67" & "1001" => d <= "11001100"; -- ##..##..
                when x"67" & "1010" => d <= "11001100"; -- ##..##..
                when x"67" & "1011" => d <= "01111100"; -- .#####..
                when x"67" & "1100" => d <= "00001100"; -- ....##..
                when x"67" & "1101" => d <= "11001100"; -- ##..##..
                when x"67" & "1110" => d <= "01111000"; -- .####...
                when x"67" & "1111" => d <= "00000000"; -- ........

                when x"68" & "0000" => d <= "00000000"; -- ........
                when x"68" & "0001" => d <= "00000000"; -- ........
                when x"68" & "0010" => d <= "11100000"; -- ###.....
                when x"68" & "0011" => d <= "01100000"; -- .##.....
                when x"68" & "0100" => d <= "01100000"; -- .##.....
                when x"68" & "0101" => d <= "01101100"; -- .##.##..
                when x"68" & "0110" => d <= "01110110"; -- .###.##.
                when x"68" & "0111" => d <= "01100110"; -- .##..##.
                when x"68" & "1000" => d <= "01100110"; -- .##..##.
                when x"68" & "1001" => d <= "01100110"; -- .##..##.
                when x"68" & "1010" => d <= "01100110"; -- .##..##.
                when x"68" & "1011" => d <= "11100110"; -- ###..##.
                when x"68" & "1100" => d <= "00000000"; -- ........
                when x"68" & "1101" => d <= "00000000"; -- ........
                when x"68" & "1110" => d <= "00000000"; -- ........
                when x"68" & "1111" => d <= "00000000"; -- ........

                when x"69" & "0000" => d <= "00000000"; -- ........
                when x"69" & "0001" => d <= "00000000"; -- ........
                when x"69" & "0010" => d <= "00011000"; -- ...##...
                when x"69" & "0011" => d <= "00011000"; -- ...##...
                when x"69" & "0100" => d <= "00000000"; -- ........
                when x"69" & "0101" => d <= "00111000"; -- ..###...
                when x"69" & "0110" => d <= "00011000"; -- ...##...
                when x"69" & "0111" => d <= "00011000"; -- ...##...
                when x"69" & "1000" => d <= "00011000"; -- ...##...
                when x"69" & "1001" => d <= "00011000"; -- ...##...
                when x"69" & "1010" => d <= "00011000"; -- ...##...
                when x"69" & "1011" => d <= "00111100"; -- ..####..
                when x"69" & "1100" => d <= "00000000"; -- ........
                when x"69" & "1101" => d <= "00000000"; -- ........
                when x"69" & "1110" => d <= "00000000"; -- ........
                when x"69" & "1111" => d <= "00000000"; -- ........

                when x"6a" & "0000" => d <= "00000000"; -- ........
                when x"6a" & "0001" => d <= "00000000"; -- ........
                when x"6a" & "0010" => d <= "00000110"; -- .....##.
                when x"6a" & "0011" => d <= "00000110"; -- .....##.
                when x"6a" & "0100" => d <= "00000000"; -- ........
                when x"6a" & "0101" => d <= "00001110"; -- ....###.
                when x"6a" & "0110" => d <= "00000110"; -- .....##.
                when x"6a" & "0111" => d <= "00000110"; -- .....##.
                when x"6a" & "1000" => d <= "00000110"; -- .....##.
                when x"6a" & "1001" => d <= "00000110"; -- .....##.
                when x"6a" & "1010" => d <= "00000110"; -- .....##.
                when x"6a" & "1011" => d <= "00000110"; -- .....##.
                when x"6a" & "1100" => d <= "01100110"; -- .##..##.
                when x"6a" & "1101" => d <= "01100110"; -- .##..##.
                when x"6a" & "1110" => d <= "00111100"; -- ..####..
                when x"6a" & "1111" => d <= "00000000"; -- ........

                when x"6b" & "0000" => d <= "00000000"; -- ........
                when x"6b" & "0001" => d <= "00000000"; -- ........
                when x"6b" & "0010" => d <= "11100000"; -- ###.....
                when x"6b" & "0011" => d <= "01100000"; -- .##.....
                when x"6b" & "0100" => d <= "01100000"; -- .##.....
                when x"6b" & "0101" => d <= "01100110"; -- .##..##.
                when x"6b" & "0110" => d <= "01101100"; -- .##.##..
                when x"6b" & "0111" => d <= "01111000"; -- .####...
                when x"6b" & "1000" => d <= "01111000"; -- .####...
                when x"6b" & "1001" => d <= "01101100"; -- .##.##..
                when x"6b" & "1010" => d <= "01100110"; -- .##..##.
                when x"6b" & "1011" => d <= "11100110"; -- ###..##.
                when x"6b" & "1100" => d <= "00000000"; -- ........
                when x"6b" & "1101" => d <= "00000000"; -- ........
                when x"6b" & "1110" => d <= "00000000"; -- ........
                when x"6b" & "1111" => d <= "00000000"; -- ........

                when x"6c" & "0000" => d <= "00000000"; -- ........
                when x"6c" & "0001" => d <= "00000000"; -- ........
                when x"6c" & "0010" => d <= "00111000"; -- ..###...
                when x"6c" & "0011" => d <= "00011000"; -- ...##...
                when x"6c" & "0100" => d <= "00011000"; -- ...##...
                when x"6c" & "0101" => d <= "00011000"; -- ...##...
                when x"6c" & "0110" => d <= "00011000"; -- ...##...
                when x"6c" & "0111" => d <= "00011000"; -- ...##...
                when x"6c" & "1000" => d <= "00011000"; -- ...##...
                when x"6c" & "1001" => d <= "00011000"; -- ...##...
                when x"6c" & "1010" => d <= "00011000"; -- ...##...
                when x"6c" & "1011" => d <= "00111100"; -- ..####..
                when x"6c" & "1100" => d <= "00000000"; -- ........
                when x"6c" & "1101" => d <= "00000000"; -- ........
                when x"6c" & "1110" => d <= "00000000"; -- ........
                when x"6c" & "1111" => d <= "00000000"; -- ........

                when x"6d" & "0000" => d <= "00000000"; -- ........
                when x"6d" & "0001" => d <= "00000000"; -- ........
                when x"6d" & "0010" => d <= "00000000"; -- ........
                when x"6d" & "0011" => d <= "00000000"; -- ........
                when x"6d" & "0100" => d <= "00000000"; -- ........
                when x"6d" & "0101" => d <= "11101100"; -- ###.##..
                when x"6d" & "0110" => d <= "11111110"; -- #######.
                when x"6d" & "0111" => d <= "11010110"; -- ##.#.##.
                when x"6d" & "1000" => d <= "11010110"; -- ##.#.##.
                when x"6d" & "1001" => d <= "11010110"; -- ##.#.##.
                when x"6d" & "1010" => d <= "11010110"; -- ##.#.##.
                when x"6d" & "1011" => d <= "11000110"; -- ##...##.
                when x"6d" & "1100" => d <= "00000000"; -- ........
                when x"6d" & "1101" => d <= "00000000"; -- ........
                when x"6d" & "1110" => d <= "00000000"; -- ........
                when x"6d" & "1111" => d <= "00000000"; -- ........

                when x"6e" & "0000" => d <= "00000000"; -- ........
                when x"6e" & "0001" => d <= "00000000"; -- ........
                when x"6e" & "0010" => d <= "00000000"; -- ........
                when x"6e" & "0011" => d <= "00000000"; -- ........
                when x"6e" & "0100" => d <= "00000000"; -- ........
                when x"6e" & "0101" => d <= "11011100"; -- ##.###..
                when x"6e" & "0110" => d <= "01100110"; -- .##..##.
                when x"6e" & "0111" => d <= "01100110"; -- .##..##.
                when x"6e" & "1000" => d <= "01100110"; -- .##..##.
                when x"6e" & "1001" => d <= "01100110"; -- .##..##.
                when x"6e" & "1010" => d <= "01100110"; -- .##..##.
                when x"6e" & "1011" => d <= "01100110"; -- .##..##.
                when x"6e" & "1100" => d <= "00000000"; -- ........
                when x"6e" & "1101" => d <= "00000000"; -- ........
                when x"6e" & "1110" => d <= "00000000"; -- ........
                when x"6e" & "1111" => d <= "00000000"; -- ........

                when x"6f" & "0000" => d <= "00000000"; -- ........
                when x"6f" & "0001" => d <= "00000000"; -- ........
                when x"6f" & "0010" => d <= "00000000"; -- ........
                when x"6f" & "0011" => d <= "00000000"; -- ........
                when x"6f" & "0100" => d <= "00000000"; -- ........
                when x"6f" & "0101" => d <= "01111100"; -- .#####..
                when x"6f" & "0110" => d <= "11000110"; -- ##...##.
                when x"6f" & "0111" => d <= "11000110"; -- ##...##.
                when x"6f" & "1000" => d <= "11000110"; -- ##...##.
                when x"6f" & "1001" => d <= "11000110"; -- ##...##.
                when x"6f" & "1010" => d <= "11000110"; -- ##...##.
                when x"6f" & "1011" => d <= "01111100"; -- .#####..
                when x"6f" & "1100" => d <= "00000000"; -- ........
                when x"6f" & "1101" => d <= "00000000"; -- ........
                when x"6f" & "1110" => d <= "00000000"; -- ........
                when x"6f" & "1111" => d <= "00000000"; -- ........

                when x"70" & "0000" => d <= "00000000"; -- ........
                when x"70" & "0001" => d <= "00000000"; -- ........
                when x"70" & "0010" => d <= "00000000"; -- ........
                when x"70" & "0011" => d <= "00000000"; -- ........
                when x"70" & "0100" => d <= "00000000"; -- ........
                when x"70" & "0101" => d <= "11011100"; -- ##.###..
                when x"70" & "0110" => d <= "01100110"; -- .##..##.
                when x"70" & "0111" => d <= "01100110"; -- .##..##.
                when x"70" & "1000" => d <= "01100110"; -- .##..##.
                when x"70" & "1001" => d <= "01100110"; -- .##..##.
                when x"70" & "1010" => d <= "01100110"; -- .##..##.
                when x"70" & "1011" => d <= "01111100"; -- .#####..
                when x"70" & "1100" => d <= "01100000"; -- .##.....
                when x"70" & "1101" => d <= "01100000"; -- .##.....
                when x"70" & "1110" => d <= "11110000"; -- ####....
                when x"70" & "1111" => d <= "00000000"; -- ........

                when x"71" & "0000" => d <= "00000000"; -- ........
                when x"71" & "0001" => d <= "00000000"; -- ........
                when x"71" & "0010" => d <= "00000000"; -- ........
                when x"71" & "0011" => d <= "00000000"; -- ........
                when x"71" & "0100" => d <= "00000000"; -- ........
                when x"71" & "0101" => d <= "01110110"; -- .###.##.
                when x"71" & "0110" => d <= "11001100"; -- ##..##..
                when x"71" & "0111" => d <= "11001100"; -- ##..##..
                when x"71" & "1000" => d <= "11001100"; -- ##..##..
                when x"71" & "1001" => d <= "11001100"; -- ##..##..
                when x"71" & "1010" => d <= "11001100"; -- ##..##..
                when x"71" & "1011" => d <= "01111100"; -- .#####..
                when x"71" & "1100" => d <= "00001100"; -- ....##..
                when x"71" & "1101" => d <= "00001100"; -- ....##..
                when x"71" & "1110" => d <= "00011110"; -- ...####.
                when x"71" & "1111" => d <= "00000000"; -- ........

                when x"72" & "0000" => d <= "00000000"; -- ........
                when x"72" & "0001" => d <= "00000000"; -- ........
                when x"72" & "0010" => d <= "00000000"; -- ........
                when x"72" & "0011" => d <= "00000000"; -- ........
                when x"72" & "0100" => d <= "00000000"; -- ........
                when x"72" & "0101" => d <= "11011100"; -- ##.###..
                when x"72" & "0110" => d <= "01110110"; -- .###.##.
                when x"72" & "0111" => d <= "01100110"; -- .##..##.
                when x"72" & "1000" => d <= "01100000"; -- .##.....
                when x"72" & "1001" => d <= "01100000"; -- .##.....
                when x"72" & "1010" => d <= "01100000"; -- .##.....
                when x"72" & "1011" => d <= "11110000"; -- ####....
                when x"72" & "1100" => d <= "00000000"; -- ........
                when x"72" & "1101" => d <= "00000000"; -- ........
                when x"72" & "1110" => d <= "00000000"; -- ........
                when x"72" & "1111" => d <= "00000000"; -- ........

                when x"73" & "0000" => d <= "00000000"; -- ........
                when x"73" & "0001" => d <= "00000000"; -- ........
                when x"73" & "0010" => d <= "00000000"; -- ........
                when x"73" & "0011" => d <= "00000000"; -- ........
                when x"73" & "0100" => d <= "00000000"; -- ........
                when x"73" & "0101" => d <= "01111100"; -- .#####..
                when x"73" & "0110" => d <= "11000110"; -- ##...##.
                when x"73" & "0111" => d <= "01100000"; -- .##.....
                when x"73" & "1000" => d <= "00111000"; -- ..###...
                when x"73" & "1001" => d <= "00001100"; -- ....##..
                when x"73" & "1010" => d <= "11000110"; -- ##...##.
                when x"73" & "1011" => d <= "01111100"; -- .#####..
                when x"73" & "1100" => d <= "00000000"; -- ........
                when x"73" & "1101" => d <= "00000000"; -- ........
                when x"73" & "1110" => d <= "00000000"; -- ........
                when x"73" & "1111" => d <= "00000000"; -- ........

                when x"74" & "0000" => d <= "00000000"; -- ........
                when x"74" & "0001" => d <= "00000000"; -- ........
                when x"74" & "0010" => d <= "00010000"; -- ...#....
                when x"74" & "0011" => d <= "00110000"; -- ..##....
                when x"74" & "0100" => d <= "00110000"; -- ..##....
                when x"74" & "0101" => d <= "11111100"; -- ######..
                when x"74" & "0110" => d <= "00110000"; -- ..##....
                when x"74" & "0111" => d <= "00110000"; -- ..##....
                when x"74" & "1000" => d <= "00110000"; -- ..##....
                when x"74" & "1001" => d <= "00110000"; -- ..##....
                when x"74" & "1010" => d <= "00110110"; -- ..##.##.
                when x"74" & "1011" => d <= "00011100"; -- ...###..
                when x"74" & "1100" => d <= "00000000"; -- ........
                when x"74" & "1101" => d <= "00000000"; -- ........
                when x"74" & "1110" => d <= "00000000"; -- ........
                when x"74" & "1111" => d <= "00000000"; -- ........

                when x"75" & "0000" => d <= "00000000"; -- ........
                when x"75" & "0001" => d <= "00000000"; -- ........
                when x"75" & "0010" => d <= "00000000"; -- ........
                when x"75" & "0011" => d <= "00000000"; -- ........
                when x"75" & "0100" => d <= "00000000"; -- ........
                when x"75" & "0101" => d <= "11001100"; -- ##..##..
                when x"75" & "0110" => d <= "11001100"; -- ##..##..
                when x"75" & "0111" => d <= "11001100"; -- ##..##..
                when x"75" & "1000" => d <= "11001100"; -- ##..##..
                when x"75" & "1001" => d <= "11001100"; -- ##..##..
                when x"75" & "1010" => d <= "11001100"; -- ##..##..
                when x"75" & "1011" => d <= "01110110"; -- .###.##.
                when x"75" & "1100" => d <= "00000000"; -- ........
                when x"75" & "1101" => d <= "00000000"; -- ........
                when x"75" & "1110" => d <= "00000000"; -- ........
                when x"75" & "1111" => d <= "00000000"; -- ........

                when x"76" & "0000" => d <= "00000000"; -- ........
                when x"76" & "0001" => d <= "00000000"; -- ........
                when x"76" & "0010" => d <= "00000000"; -- ........
                when x"76" & "0011" => d <= "00000000"; -- ........
                when x"76" & "0100" => d <= "00000000"; -- ........
                when x"76" & "0101" => d <= "01100110"; -- .##..##.
                when x"76" & "0110" => d <= "01100110"; -- .##..##.
                when x"76" & "0111" => d <= "01100110"; -- .##..##.
                when x"76" & "1000" => d <= "01100110"; -- .##..##.
                when x"76" & "1001" => d <= "01100110"; -- .##..##.
                when x"76" & "1010" => d <= "00111100"; -- ..####..
                when x"76" & "1011" => d <= "00011000"; -- ...##...
                when x"76" & "1100" => d <= "00000000"; -- ........
                when x"76" & "1101" => d <= "00000000"; -- ........
                when x"76" & "1110" => d <= "00000000"; -- ........
                when x"76" & "1111" => d <= "00000000"; -- ........

                when x"77" & "0000" => d <= "00000000"; -- ........
                when x"77" & "0001" => d <= "00000000"; -- ........
                when x"77" & "0010" => d <= "00000000"; -- ........
                when x"77" & "0011" => d <= "00000000"; -- ........
                when x"77" & "0100" => d <= "00000000"; -- ........
                when x"77" & "0101" => d <= "11000110"; -- ##...##.
                when x"77" & "0110" => d <= "11000110"; -- ##...##.
                when x"77" & "0111" => d <= "11010110"; -- ##.#.##.
                when x"77" & "1000" => d <= "11010110"; -- ##.#.##.
                when x"77" & "1001" => d <= "11010110"; -- ##.#.##.
                when x"77" & "1010" => d <= "11111110"; -- #######.
                when x"77" & "1011" => d <= "01101100"; -- .##.##..
                when x"77" & "1100" => d <= "00000000"; -- ........
                when x"77" & "1101" => d <= "00000000"; -- ........
                when x"77" & "1110" => d <= "00000000"; -- ........
                when x"77" & "1111" => d <= "00000000"; -- ........

                when x"78" & "0000" => d <= "00000000"; -- ........
                when x"78" & "0001" => d <= "00000000"; -- ........
                when x"78" & "0010" => d <= "00000000"; -- ........
                when x"78" & "0011" => d <= "00000000"; -- ........
                when x"78" & "0100" => d <= "00000000"; -- ........
                when x"78" & "0101" => d <= "11000110"; -- ##...##.
                when x"78" & "0110" => d <= "01101100"; -- .##.##..
                when x"78" & "0111" => d <= "00111000"; -- ..###...
                when x"78" & "1000" => d <= "00111000"; -- ..###...
                when x"78" & "1001" => d <= "00111000"; -- ..###...
                when x"78" & "1010" => d <= "01101100"; -- .##.##..
                when x"78" & "1011" => d <= "11000110"; -- ##...##.
                when x"78" & "1100" => d <= "00000000"; -- ........
                when x"78" & "1101" => d <= "00000000"; -- ........
                when x"78" & "1110" => d <= "00000000"; -- ........
                when x"78" & "1111" => d <= "00000000"; -- ........

                when x"79" & "0000" => d <= "00000000"; -- ........
                when x"79" & "0001" => d <= "00000000"; -- ........
                when x"79" & "0010" => d <= "00000000"; -- ........
                when x"79" & "0011" => d <= "00000000"; -- ........
                when x"79" & "0100" => d <= "00000000"; -- ........
                when x"79" & "0101" => d <= "11000110"; -- ##...##.
                when x"79" & "0110" => d <= "11000110"; -- ##...##.
                when x"79" & "0111" => d <= "11000110"; -- ##...##.
                when x"79" & "1000" => d <= "11000110"; -- ##...##.
                when x"79" & "1001" => d <= "11000110"; -- ##...##.
                when x"79" & "1010" => d <= "11000110"; -- ##...##.
                when x"79" & "1011" => d <= "01111110"; -- .######.
                when x"79" & "1100" => d <= "00000110"; -- .....##.
                when x"79" & "1101" => d <= "00001100"; -- ....##..
                when x"79" & "1110" => d <= "11111000"; -- #####...
                when x"79" & "1111" => d <= "00000000"; -- ........

                when x"7a" & "0000" => d <= "00000000"; -- ........
                when x"7a" & "0001" => d <= "00000000"; -- ........
                when x"7a" & "0010" => d <= "00000000"; -- ........
                when x"7a" & "0011" => d <= "00000000"; -- ........
                when x"7a" & "0100" => d <= "00000000"; -- ........
                when x"7a" & "0101" => d <= "11111110"; -- #######.
                when x"7a" & "0110" => d <= "11001100"; -- ##..##..
                when x"7a" & "0111" => d <= "00011000"; -- ...##...
                when x"7a" & "1000" => d <= "00110000"; -- ..##....
                when x"7a" & "1001" => d <= "01100000"; -- .##.....
                when x"7a" & "1010" => d <= "11000110"; -- ##...##.
                when x"7a" & "1011" => d <= "11111110"; -- #######.
                when x"7a" & "1100" => d <= "00000000"; -- ........
                when x"7a" & "1101" => d <= "00000000"; -- ........
                when x"7a" & "1110" => d <= "00000000"; -- ........
                when x"7a" & "1111" => d <= "00000000"; -- ........

                when x"7b" & "0000" => d <= "00000000"; -- ........
                when x"7b" & "0001" => d <= "00000000"; -- ........
                when x"7b" & "0010" => d <= "00001110"; -- ....###.
                when x"7b" & "0011" => d <= "00011000"; -- ...##...
                when x"7b" & "0100" => d <= "00011000"; -- ...##...
                when x"7b" & "0101" => d <= "00011000"; -- ...##...
                when x"7b" & "0110" => d <= "01110000"; -- .###....
                when x"7b" & "0111" => d <= "00011000"; -- ...##...
                when x"7b" & "1000" => d <= "00011000"; -- ...##...
                when x"7b" & "1001" => d <= "00011000"; -- ...##...
                when x"7b" & "1010" => d <= "00011000"; -- ...##...
                when x"7b" & "1011" => d <= "00001110"; -- ....###.
                when x"7b" & "1100" => d <= "00000000"; -- ........
                when x"7b" & "1101" => d <= "00000000"; -- ........
                when x"7b" & "1110" => d <= "00000000"; -- ........
                when x"7b" & "1111" => d <= "00000000"; -- ........

                when x"7c" & "0000" => d <= "00000000"; -- ........
                when x"7c" & "0001" => d <= "00000000"; -- ........
                when x"7c" & "0010" => d <= "00011000"; -- ...##...
                when x"7c" & "0011" => d <= "00011000"; -- ...##...
                when x"7c" & "0100" => d <= "00011000"; -- ...##...
                when x"7c" & "0101" => d <= "00011000"; -- ...##...
                when x"7c" & "0110" => d <= "00000000"; -- ........
                when x"7c" & "0111" => d <= "00011000"; -- ...##...
                when x"7c" & "1000" => d <= "00011000"; -- ...##...
                when x"7c" & "1001" => d <= "00011000"; -- ...##...
                when x"7c" & "1010" => d <= "00011000"; -- ...##...
                when x"7c" & "1011" => d <= "00011000"; -- ...##...
                when x"7c" & "1100" => d <= "00000000"; -- ........
                when x"7c" & "1101" => d <= "00000000"; -- ........
                when x"7c" & "1110" => d <= "00000000"; -- ........
                when x"7c" & "1111" => d <= "00000000"; -- ........

                when x"7d" & "0000" => d <= "00000000"; -- ........
                when x"7d" & "0001" => d <= "00000000"; -- ........
                when x"7d" & "0010" => d <= "01110000"; -- .###....
                when x"7d" & "0011" => d <= "00011000"; -- ...##...
                when x"7d" & "0100" => d <= "00011000"; -- ...##...
                when x"7d" & "0101" => d <= "00011000"; -- ...##...
                when x"7d" & "0110" => d <= "00001110"; -- ....###.
                when x"7d" & "0111" => d <= "00011000"; -- ...##...
                when x"7d" & "1000" => d <= "00011000"; -- ...##...
                when x"7d" & "1001" => d <= "00011000"; -- ...##...
                when x"7d" & "1010" => d <= "00011000"; -- ...##...
                when x"7d" & "1011" => d <= "01110000"; -- .###....
                when x"7d" & "1100" => d <= "00000000"; -- ........
                when x"7d" & "1101" => d <= "00000000"; -- ........
                when x"7d" & "1110" => d <= "00000000"; -- ........
                when x"7d" & "1111" => d <= "00000000"; -- ........

                when x"7e" & "0000" => d <= "00000000"; -- ........
                when x"7e" & "0001" => d <= "00000000"; -- ........
                when x"7e" & "0010" => d <= "01110110"; -- .###.##.
                when x"7e" & "0011" => d <= "11011100"; -- ##.###..
                when x"7e" & "0100" => d <= "00000000"; -- ........
                when x"7e" & "0101" => d <= "00000000"; -- ........
                when x"7e" & "0110" => d <= "00000000"; -- ........
                when x"7e" & "0111" => d <= "00000000"; -- ........
                when x"7e" & "1000" => d <= "00000000"; -- ........
                when x"7e" & "1001" => d <= "00000000"; -- ........
                when x"7e" & "1010" => d <= "00000000"; -- ........
                when x"7e" & "1011" => d <= "00000000"; -- ........
                when x"7e" & "1100" => d <= "00000000"; -- ........
                when x"7e" & "1101" => d <= "00000000"; -- ........
                when x"7e" & "1110" => d <= "00000000"; -- ........
                when x"7e" & "1111" => d <= "00000000"; -- ........

                when x"7f" & "0000" => d <= "00000000"; -- ........
                when x"7f" & "0001" => d <= "00000000"; -- ........
                when x"7f" & "0010" => d <= "00000000"; -- ........
                when x"7f" & "0011" => d <= "00000000"; -- ........
                when x"7f" & "0100" => d <= "00010000"; -- ...#....
                when x"7f" & "0101" => d <= "00111000"; -- ..###...
                when x"7f" & "0110" => d <= "01101100"; -- .##.##..
                when x"7f" & "0111" => d <= "11000110"; -- ##...##.
                when x"7f" & "1000" => d <= "11000110"; -- ##...##.
                when x"7f" & "1001" => d <= "11000110"; -- ##...##.
                when x"7f" & "1010" => d <= "11111110"; -- #######.
                when x"7f" & "1011" => d <= "00000000"; -- ........
                when x"7f" & "1100" => d <= "00000000"; -- ........
                when x"7f" & "1101" => d <= "00000000"; -- ........
                when x"7f" & "1110" => d <= "00000000"; -- ........
                when x"7f" & "1111" => d <= "00000000"; -- ........

                when x"80" & "0000" => d <= "00000000"; -- ........
                when x"80" & "0001" => d <= "00000000"; -- ........
                when x"80" & "0010" => d <= "00111100"; -- ..####..
                when x"80" & "0011" => d <= "01100110"; -- .##..##.
                when x"80" & "0100" => d <= "11000010"; -- ##....#.
                when x"80" & "0101" => d <= "11000000"; -- ##......
                when x"80" & "0110" => d <= "11000000"; -- ##......
                when x"80" & "0111" => d <= "11000000"; -- ##......
                when x"80" & "1000" => d <= "11000010"; -- ##....#.
                when x"80" & "1001" => d <= "01100110"; -- .##..##.
                when x"80" & "1010" => d <= "00111100"; -- ..####..
                when x"80" & "1011" => d <= "00001100"; -- ....##..
                when x"80" & "1100" => d <= "00000110"; -- .....##.
                when x"80" & "1101" => d <= "01111100"; -- .#####..
                when x"80" & "1110" => d <= "00000000"; -- ........
                when x"80" & "1111" => d <= "00000000"; -- ........

                when x"81" & "0000" => d <= "00000000"; -- ........
                when x"81" & "0001" => d <= "00000000"; -- ........
                when x"81" & "0010" => d <= "11001100"; -- ##..##..
                when x"81" & "0011" => d <= "00000000"; -- ........
                when x"81" & "0100" => d <= "00000000"; -- ........
                when x"81" & "0101" => d <= "11001100"; -- ##..##..
                when x"81" & "0110" => d <= "11001100"; -- ##..##..
                when x"81" & "0111" => d <= "11001100"; -- ##..##..
                when x"81" & "1000" => d <= "11001100"; -- ##..##..
                when x"81" & "1001" => d <= "11001100"; -- ##..##..
                when x"81" & "1010" => d <= "11001100"; -- ##..##..
                when x"81" & "1011" => d <= "01110110"; -- .###.##.
                when x"81" & "1100" => d <= "00000000"; -- ........
                when x"81" & "1101" => d <= "00000000"; -- ........
                when x"81" & "1110" => d <= "00000000"; -- ........
                when x"81" & "1111" => d <= "00000000"; -- ........

                when x"82" & "0000" => d <= "00000000"; -- ........
                when x"82" & "0001" => d <= "00001100"; -- ....##..
                when x"82" & "0010" => d <= "00011000"; -- ...##...
                when x"82" & "0011" => d <= "00110000"; -- ..##....
                when x"82" & "0100" => d <= "00000000"; -- ........
                when x"82" & "0101" => d <= "01111100"; -- .#####..
                when x"82" & "0110" => d <= "11000110"; -- ##...##.
                when x"82" & "0111" => d <= "11111110"; -- #######.
                when x"82" & "1000" => d <= "11000000"; -- ##......
                when x"82" & "1001" => d <= "11000000"; -- ##......
                when x"82" & "1010" => d <= "11000110"; -- ##...##.
                when x"82" & "1011" => d <= "01111100"; -- .#####..
                when x"82" & "1100" => d <= "00000000"; -- ........
                when x"82" & "1101" => d <= "00000000"; -- ........
                when x"82" & "1110" => d <= "00000000"; -- ........
                when x"82" & "1111" => d <= "00000000"; -- ........

                when x"83" & "0000" => d <= "00000000"; -- ........
                when x"83" & "0001" => d <= "00010000"; -- ...#....
                when x"83" & "0010" => d <= "00111000"; -- ..###...
                when x"83" & "0011" => d <= "01101100"; -- .##.##..
                when x"83" & "0100" => d <= "00000000"; -- ........
                when x"83" & "0101" => d <= "01111000"; -- .####...
                when x"83" & "0110" => d <= "00001100"; -- ....##..
                when x"83" & "0111" => d <= "01111100"; -- .#####..
                when x"83" & "1000" => d <= "11001100"; -- ##..##..
                when x"83" & "1001" => d <= "11001100"; -- ##..##..
                when x"83" & "1010" => d <= "11001100"; -- ##..##..
                when x"83" & "1011" => d <= "01110110"; -- .###.##.
                when x"83" & "1100" => d <= "00000000"; -- ........
                when x"83" & "1101" => d <= "00000000"; -- ........
                when x"83" & "1110" => d <= "00000000"; -- ........
                when x"83" & "1111" => d <= "00000000"; -- ........

                when x"84" & "0000" => d <= "00000000"; -- ........
                when x"84" & "0001" => d <= "00000000"; -- ........
                when x"84" & "0010" => d <= "11001100"; -- ##..##..
                when x"84" & "0011" => d <= "00000000"; -- ........
                when x"84" & "0100" => d <= "00000000"; -- ........
                when x"84" & "0101" => d <= "01111000"; -- .####...
                when x"84" & "0110" => d <= "00001100"; -- ....##..
                when x"84" & "0111" => d <= "01111100"; -- .#####..
                when x"84" & "1000" => d <= "11001100"; -- ##..##..
                when x"84" & "1001" => d <= "11001100"; -- ##..##..
                when x"84" & "1010" => d <= "11001100"; -- ##..##..
                when x"84" & "1011" => d <= "01110110"; -- .###.##.
                when x"84" & "1100" => d <= "00000000"; -- ........
                when x"84" & "1101" => d <= "00000000"; -- ........
                when x"84" & "1110" => d <= "00000000"; -- ........
                when x"84" & "1111" => d <= "00000000"; -- ........

                when x"85" & "0000" => d <= "00000000"; -- ........
                when x"85" & "0001" => d <= "01100000"; -- .##.....
                when x"85" & "0010" => d <= "00110000"; -- ..##....
                when x"85" & "0011" => d <= "00011000"; -- ...##...
                when x"85" & "0100" => d <= "00000000"; -- ........
                when x"85" & "0101" => d <= "01111000"; -- .####...
                when x"85" & "0110" => d <= "00001100"; -- ....##..
                when x"85" & "0111" => d <= "01111100"; -- .#####..
                when x"85" & "1000" => d <= "11001100"; -- ##..##..
                when x"85" & "1001" => d <= "11001100"; -- ##..##..
                when x"85" & "1010" => d <= "11001100"; -- ##..##..
                when x"85" & "1011" => d <= "01110110"; -- .###.##.
                when x"85" & "1100" => d <= "00000000"; -- ........
                when x"85" & "1101" => d <= "00000000"; -- ........
                when x"85" & "1110" => d <= "00000000"; -- ........
                when x"85" & "1111" => d <= "00000000"; -- ........

                when x"86" & "0000" => d <= "00000000"; -- ........
                when x"86" & "0001" => d <= "00111000"; -- ..###...
                when x"86" & "0010" => d <= "01101100"; -- .##.##..
                when x"86" & "0011" => d <= "00111000"; -- ..###...
                when x"86" & "0100" => d <= "00000000"; -- ........
                when x"86" & "0101" => d <= "01111000"; -- .####...
                when x"86" & "0110" => d <= "00001100"; -- ....##..
                when x"86" & "0111" => d <= "01111100"; -- .#####..
                when x"86" & "1000" => d <= "11001100"; -- ##..##..
                when x"86" & "1001" => d <= "11001100"; -- ##..##..
                when x"86" & "1010" => d <= "11001100"; -- ##..##..
                when x"86" & "1011" => d <= "01110110"; -- .###.##.
                when x"86" & "1100" => d <= "00000000"; -- ........
                when x"86" & "1101" => d <= "00000000"; -- ........
                when x"86" & "1110" => d <= "00000000"; -- ........
                when x"86" & "1111" => d <= "00000000"; -- ........

                when x"87" & "0000" => d <= "00000000"; -- ........
                when x"87" & "0001" => d <= "00000000"; -- ........
                when x"87" & "0010" => d <= "00000000"; -- ........
                when x"87" & "0011" => d <= "00000000"; -- ........
                when x"87" & "0100" => d <= "00111100"; -- ..####..
                when x"87" & "0101" => d <= "01100110"; -- .##..##.
                when x"87" & "0110" => d <= "01100000"; -- .##.....
                when x"87" & "0111" => d <= "01100000"; -- .##.....
                when x"87" & "1000" => d <= "01100110"; -- .##..##.
                when x"87" & "1001" => d <= "00111100"; -- ..####..
                when x"87" & "1010" => d <= "00001100"; -- ....##..
                when x"87" & "1011" => d <= "00000110"; -- .....##.
                when x"87" & "1100" => d <= "00111100"; -- ..####..
                when x"87" & "1101" => d <= "00000000"; -- ........
                when x"87" & "1110" => d <= "00000000"; -- ........
                when x"87" & "1111" => d <= "00000000"; -- ........

                when x"88" & "0000" => d <= "00000000"; -- ........
                when x"88" & "0001" => d <= "00010000"; -- ...#....
                when x"88" & "0010" => d <= "00111000"; -- ..###...
                when x"88" & "0011" => d <= "01101100"; -- .##.##..
                when x"88" & "0100" => d <= "00000000"; -- ........
                when x"88" & "0101" => d <= "01111100"; -- .#####..
                when x"88" & "0110" => d <= "11000110"; -- ##...##.
                when x"88" & "0111" => d <= "11111110"; -- #######.
                when x"88" & "1000" => d <= "11000000"; -- ##......
                when x"88" & "1001" => d <= "11000000"; -- ##......
                when x"88" & "1010" => d <= "11000110"; -- ##...##.
                when x"88" & "1011" => d <= "01111100"; -- .#####..
                when x"88" & "1100" => d <= "00000000"; -- ........
                when x"88" & "1101" => d <= "00000000"; -- ........
                when x"88" & "1110" => d <= "00000000"; -- ........
                when x"88" & "1111" => d <= "00000000"; -- ........

                when x"89" & "0000" => d <= "00000000"; -- ........
                when x"89" & "0001" => d <= "00000000"; -- ........
                when x"89" & "0010" => d <= "11000110"; -- ##...##.
                when x"89" & "0011" => d <= "00000000"; -- ........
                when x"89" & "0100" => d <= "00000000"; -- ........
                when x"89" & "0101" => d <= "01111100"; -- .#####..
                when x"89" & "0110" => d <= "11000110"; -- ##...##.
                when x"89" & "0111" => d <= "11111110"; -- #######.
                when x"89" & "1000" => d <= "11000000"; -- ##......
                when x"89" & "1001" => d <= "11000000"; -- ##......
                when x"89" & "1010" => d <= "11000110"; -- ##...##.
                when x"89" & "1011" => d <= "01111100"; -- .#####..
                when x"89" & "1100" => d <= "00000000"; -- ........
                when x"89" & "1101" => d <= "00000000"; -- ........
                when x"89" & "1110" => d <= "00000000"; -- ........
                when x"89" & "1111" => d <= "00000000"; -- ........

                when x"8a" & "0000" => d <= "00000000"; -- ........
                when x"8a" & "0001" => d <= "01100000"; -- .##.....
                when x"8a" & "0010" => d <= "00110000"; -- ..##....
                when x"8a" & "0011" => d <= "00011000"; -- ...##...
                when x"8a" & "0100" => d <= "00000000"; -- ........
                when x"8a" & "0101" => d <= "01111100"; -- .#####..
                when x"8a" & "0110" => d <= "11000110"; -- ##...##.
                when x"8a" & "0111" => d <= "11111110"; -- #######.
                when x"8a" & "1000" => d <= "11000000"; -- ##......
                when x"8a" & "1001" => d <= "11000000"; -- ##......
                when x"8a" & "1010" => d <= "11000110"; -- ##...##.
                when x"8a" & "1011" => d <= "01111100"; -- .#####..
                when x"8a" & "1100" => d <= "00000000"; -- ........
                when x"8a" & "1101" => d <= "00000000"; -- ........
                when x"8a" & "1110" => d <= "00000000"; -- ........
                when x"8a" & "1111" => d <= "00000000"; -- ........

                when x"8b" & "0000" => d <= "00000000"; -- ........
                when x"8b" & "0001" => d <= "00000000"; -- ........
                when x"8b" & "0010" => d <= "01100110"; -- .##..##.
                when x"8b" & "0011" => d <= "00000000"; -- ........
                when x"8b" & "0100" => d <= "00000000"; -- ........
                when x"8b" & "0101" => d <= "00111000"; -- ..###...
                when x"8b" & "0110" => d <= "00011000"; -- ...##...
                when x"8b" & "0111" => d <= "00011000"; -- ...##...
                when x"8b" & "1000" => d <= "00011000"; -- ...##...
                when x"8b" & "1001" => d <= "00011000"; -- ...##...
                when x"8b" & "1010" => d <= "00011000"; -- ...##...
                when x"8b" & "1011" => d <= "00111100"; -- ..####..
                when x"8b" & "1100" => d <= "00000000"; -- ........
                when x"8b" & "1101" => d <= "00000000"; -- ........
                when x"8b" & "1110" => d <= "00000000"; -- ........
                when x"8b" & "1111" => d <= "00000000"; -- ........

                when x"8c" & "0000" => d <= "00000000"; -- ........
                when x"8c" & "0001" => d <= "00011000"; -- ...##...
                when x"8c" & "0010" => d <= "00111100"; -- ..####..
                when x"8c" & "0011" => d <= "01100110"; -- .##..##.
                when x"8c" & "0100" => d <= "00000000"; -- ........
                when x"8c" & "0101" => d <= "00111000"; -- ..###...
                when x"8c" & "0110" => d <= "00011000"; -- ...##...
                when x"8c" & "0111" => d <= "00011000"; -- ...##...
                when x"8c" & "1000" => d <= "00011000"; -- ...##...
                when x"8c" & "1001" => d <= "00011000"; -- ...##...
                when x"8c" & "1010" => d <= "00011000"; -- ...##...
                when x"8c" & "1011" => d <= "00111100"; -- ..####..
                when x"8c" & "1100" => d <= "00000000"; -- ........
                when x"8c" & "1101" => d <= "00000000"; -- ........
                when x"8c" & "1110" => d <= "00000000"; -- ........
                when x"8c" & "1111" => d <= "00000000"; -- ........

                when x"8d" & "0000" => d <= "00000000"; -- ........
                when x"8d" & "0001" => d <= "01100000"; -- .##.....
                when x"8d" & "0010" => d <= "00110000"; -- ..##....
                when x"8d" & "0011" => d <= "00011000"; -- ...##...
                when x"8d" & "0100" => d <= "00000000"; -- ........
                when x"8d" & "0101" => d <= "00111000"; -- ..###...
                when x"8d" & "0110" => d <= "00011000"; -- ...##...
                when x"8d" & "0111" => d <= "00011000"; -- ...##...
                when x"8d" & "1000" => d <= "00011000"; -- ...##...
                when x"8d" & "1001" => d <= "00011000"; -- ...##...
                when x"8d" & "1010" => d <= "00011000"; -- ...##...
                when x"8d" & "1011" => d <= "00111100"; -- ..####..
                when x"8d" & "1100" => d <= "00000000"; -- ........
                when x"8d" & "1101" => d <= "00000000"; -- ........
                when x"8d" & "1110" => d <= "00000000"; -- ........
                when x"8d" & "1111" => d <= "00000000"; -- ........

                when x"8e" & "0000" => d <= "00000000"; -- ........
                when x"8e" & "0001" => d <= "11000110"; -- ##...##.
                when x"8e" & "0010" => d <= "00000000"; -- ........
                when x"8e" & "0011" => d <= "00010000"; -- ...#....
                when x"8e" & "0100" => d <= "00111000"; -- ..###...
                when x"8e" & "0101" => d <= "01101100"; -- .##.##..
                when x"8e" & "0110" => d <= "11000110"; -- ##...##.
                when x"8e" & "0111" => d <= "11000110"; -- ##...##.
                when x"8e" & "1000" => d <= "11111110"; -- #######.
                when x"8e" & "1001" => d <= "11000110"; -- ##...##.
                when x"8e" & "1010" => d <= "11000110"; -- ##...##.
                when x"8e" & "1011" => d <= "11000110"; -- ##...##.
                when x"8e" & "1100" => d <= "00000000"; -- ........
                when x"8e" & "1101" => d <= "00000000"; -- ........
                when x"8e" & "1110" => d <= "00000000"; -- ........
                when x"8e" & "1111" => d <= "00000000"; -- ........

                when x"8f" & "0000" => d <= "00111000"; -- ..###...
                when x"8f" & "0001" => d <= "01101100"; -- .##.##..
                when x"8f" & "0010" => d <= "00111000"; -- ..###...
                when x"8f" & "0011" => d <= "00000000"; -- ........
                when x"8f" & "0100" => d <= "00111000"; -- ..###...
                when x"8f" & "0101" => d <= "01101100"; -- .##.##..
                when x"8f" & "0110" => d <= "11000110"; -- ##...##.
                when x"8f" & "0111" => d <= "11000110"; -- ##...##.
                when x"8f" & "1000" => d <= "11111110"; -- #######.
                when x"8f" & "1001" => d <= "11000110"; -- ##...##.
                when x"8f" & "1010" => d <= "11000110"; -- ##...##.
                when x"8f" & "1011" => d <= "11000110"; -- ##...##.
                when x"8f" & "1100" => d <= "00000000"; -- ........
                when x"8f" & "1101" => d <= "00000000"; -- ........
                when x"8f" & "1110" => d <= "00000000"; -- ........
                when x"8f" & "1111" => d <= "00000000"; -- ........

                when x"90" & "0000" => d <= "00011000"; -- ...##...
                when x"90" & "0001" => d <= "00110000"; -- ..##....
                when x"90" & "0010" => d <= "01100000"; -- .##.....
                when x"90" & "0011" => d <= "00000000"; -- ........
                when x"90" & "0100" => d <= "11111110"; -- #######.
                when x"90" & "0101" => d <= "01100110"; -- .##..##.
                when x"90" & "0110" => d <= "01100000"; -- .##.....
                when x"90" & "0111" => d <= "01111100"; -- .#####..
                when x"90" & "1000" => d <= "01100000"; -- .##.....
                when x"90" & "1001" => d <= "01100000"; -- .##.....
                when x"90" & "1010" => d <= "01100110"; -- .##..##.
                when x"90" & "1011" => d <= "11111110"; -- #######.
                when x"90" & "1100" => d <= "00000000"; -- ........
                when x"90" & "1101" => d <= "00000000"; -- ........
                when x"90" & "1110" => d <= "00000000"; -- ........
                when x"90" & "1111" => d <= "00000000"; -- ........

                when x"91" & "0000" => d <= "00000000"; -- ........
                when x"91" & "0001" => d <= "00000000"; -- ........
                when x"91" & "0010" => d <= "00000000"; -- ........
                when x"91" & "0011" => d <= "00000000"; -- ........
                when x"91" & "0100" => d <= "00000000"; -- ........
                when x"91" & "0101" => d <= "11001100"; -- ##..##..
                when x"91" & "0110" => d <= "01110110"; -- .###.##.
                when x"91" & "0111" => d <= "00110110"; -- ..##.##.
                when x"91" & "1000" => d <= "01111110"; -- .######.
                when x"91" & "1001" => d <= "11011000"; -- ##.##...
                when x"91" & "1010" => d <= "11011000"; -- ##.##...
                when x"91" & "1011" => d <= "01101110"; -- .##.###.
                when x"91" & "1100" => d <= "00000000"; -- ........
                when x"91" & "1101" => d <= "00000000"; -- ........
                when x"91" & "1110" => d <= "00000000"; -- ........
                when x"91" & "1111" => d <= "00000000"; -- ........

                when x"92" & "0000" => d <= "00000000"; -- ........
                when x"92" & "0001" => d <= "00000000"; -- ........
                when x"92" & "0010" => d <= "00111110"; -- ..#####.
                when x"92" & "0011" => d <= "01101100"; -- .##.##..
                when x"92" & "0100" => d <= "11001100"; -- ##..##..
                when x"92" & "0101" => d <= "11001100"; -- ##..##..
                when x"92" & "0110" => d <= "11111110"; -- #######.
                when x"92" & "0111" => d <= "11001100"; -- ##..##..
                when x"92" & "1000" => d <= "11001100"; -- ##..##..
                when x"92" & "1001" => d <= "11001100"; -- ##..##..
                when x"92" & "1010" => d <= "11001100"; -- ##..##..
                when x"92" & "1011" => d <= "11001110"; -- ##..###.
                when x"92" & "1100" => d <= "00000000"; -- ........
                when x"92" & "1101" => d <= "00000000"; -- ........
                when x"92" & "1110" => d <= "00000000"; -- ........
                when x"92" & "1111" => d <= "00000000"; -- ........

                when x"93" & "0000" => d <= "00000000"; -- ........
                when x"93" & "0001" => d <= "00010000"; -- ...#....
                when x"93" & "0010" => d <= "00111000"; -- ..###...
                when x"93" & "0011" => d <= "01101100"; -- .##.##..
                when x"93" & "0100" => d <= "00000000"; -- ........
                when x"93" & "0101" => d <= "01111100"; -- .#####..
                when x"93" & "0110" => d <= "11000110"; -- ##...##.
                when x"93" & "0111" => d <= "11000110"; -- ##...##.
                when x"93" & "1000" => d <= "11000110"; -- ##...##.
                when x"93" & "1001" => d <= "11000110"; -- ##...##.
                when x"93" & "1010" => d <= "11000110"; -- ##...##.
                when x"93" & "1011" => d <= "01111100"; -- .#####..
                when x"93" & "1100" => d <= "00000000"; -- ........
                when x"93" & "1101" => d <= "00000000"; -- ........
                when x"93" & "1110" => d <= "00000000"; -- ........
                when x"93" & "1111" => d <= "00000000"; -- ........

                when x"94" & "0000" => d <= "00000000"; -- ........
                when x"94" & "0001" => d <= "00000000"; -- ........
                when x"94" & "0010" => d <= "11000110"; -- ##...##.
                when x"94" & "0011" => d <= "00000000"; -- ........
                when x"94" & "0100" => d <= "00000000"; -- ........
                when x"94" & "0101" => d <= "01111100"; -- .#####..
                when x"94" & "0110" => d <= "11000110"; -- ##...##.
                when x"94" & "0111" => d <= "11000110"; -- ##...##.
                when x"94" & "1000" => d <= "11000110"; -- ##...##.
                when x"94" & "1001" => d <= "11000110"; -- ##...##.
                when x"94" & "1010" => d <= "11000110"; -- ##...##.
                when x"94" & "1011" => d <= "01111100"; -- .#####..
                when x"94" & "1100" => d <= "00000000"; -- ........
                when x"94" & "1101" => d <= "00000000"; -- ........
                when x"94" & "1110" => d <= "00000000"; -- ........
                when x"94" & "1111" => d <= "00000000"; -- ........

                when x"95" & "0000" => d <= "00000000"; -- ........
                when x"95" & "0001" => d <= "01100000"; -- .##.....
                when x"95" & "0010" => d <= "00110000"; -- ..##....
                when x"95" & "0011" => d <= "00011000"; -- ...##...
                when x"95" & "0100" => d <= "00000000"; -- ........
                when x"95" & "0101" => d <= "01111100"; -- .#####..
                when x"95" & "0110" => d <= "11000110"; -- ##...##.
                when x"95" & "0111" => d <= "11000110"; -- ##...##.
                when x"95" & "1000" => d <= "11000110"; -- ##...##.
                when x"95" & "1001" => d <= "11000110"; -- ##...##.
                when x"95" & "1010" => d <= "11000110"; -- ##...##.
                when x"95" & "1011" => d <= "01111100"; -- .#####..
                when x"95" & "1100" => d <= "00000000"; -- ........
                when x"95" & "1101" => d <= "00000000"; -- ........
                when x"95" & "1110" => d <= "00000000"; -- ........
                when x"95" & "1111" => d <= "00000000"; -- ........

                when x"96" & "0000" => d <= "00000000"; -- ........
                when x"96" & "0001" => d <= "00110000"; -- ..##....
                when x"96" & "0010" => d <= "01111000"; -- .####...
                when x"96" & "0011" => d <= "11001100"; -- ##..##..
                when x"96" & "0100" => d <= "00000000"; -- ........
                when x"96" & "0101" => d <= "11001100"; -- ##..##..
                when x"96" & "0110" => d <= "11001100"; -- ##..##..
                when x"96" & "0111" => d <= "11001100"; -- ##..##..
                when x"96" & "1000" => d <= "11001100"; -- ##..##..
                when x"96" & "1001" => d <= "11001100"; -- ##..##..
                when x"96" & "1010" => d <= "11001100"; -- ##..##..
                when x"96" & "1011" => d <= "01110110"; -- .###.##.
                when x"96" & "1100" => d <= "00000000"; -- ........
                when x"96" & "1101" => d <= "00000000"; -- ........
                when x"96" & "1110" => d <= "00000000"; -- ........
                when x"96" & "1111" => d <= "00000000"; -- ........

                when x"97" & "0000" => d <= "00000000"; -- ........
                when x"97" & "0001" => d <= "01100000"; -- .##.....
                when x"97" & "0010" => d <= "00110000"; -- ..##....
                when x"97" & "0011" => d <= "00011000"; -- ...##...
                when x"97" & "0100" => d <= "00000000"; -- ........
                when x"97" & "0101" => d <= "11001100"; -- ##..##..
                when x"97" & "0110" => d <= "11001100"; -- ##..##..
                when x"97" & "0111" => d <= "11001100"; -- ##..##..
                when x"97" & "1000" => d <= "11001100"; -- ##..##..
                when x"97" & "1001" => d <= "11001100"; -- ##..##..
                when x"97" & "1010" => d <= "11001100"; -- ##..##..
                when x"97" & "1011" => d <= "01110110"; -- .###.##.
                when x"97" & "1100" => d <= "00000000"; -- ........
                when x"97" & "1101" => d <= "00000000"; -- ........
                when x"97" & "1110" => d <= "00000000"; -- ........
                when x"97" & "1111" => d <= "00000000"; -- ........

                when x"98" & "0000" => d <= "00000000"; -- ........
                when x"98" & "0001" => d <= "00000000"; -- ........
                when x"98" & "0010" => d <= "11000110"; -- ##...##.
                when x"98" & "0011" => d <= "00000000"; -- ........
                when x"98" & "0100" => d <= "00000000"; -- ........
                when x"98" & "0101" => d <= "11000110"; -- ##...##.
                when x"98" & "0110" => d <= "11000110"; -- ##...##.
                when x"98" & "0111" => d <= "11000110"; -- ##...##.
                when x"98" & "1000" => d <= "11000110"; -- ##...##.
                when x"98" & "1001" => d <= "11000110"; -- ##...##.
                when x"98" & "1010" => d <= "11000110"; -- ##...##.
                when x"98" & "1011" => d <= "01111110"; -- .######.
                when x"98" & "1100" => d <= "00000110"; -- .....##.
                when x"98" & "1101" => d <= "00001100"; -- ....##..
                when x"98" & "1110" => d <= "01111000"; -- .####...
                when x"98" & "1111" => d <= "00000000"; -- ........

                when x"99" & "0000" => d <= "00000000"; -- ........
                when x"99" & "0001" => d <= "11000110"; -- ##...##.
                when x"99" & "0010" => d <= "00000000"; -- ........
                when x"99" & "0011" => d <= "01111100"; -- .#####..
                when x"99" & "0100" => d <= "11000110"; -- ##...##.
                when x"99" & "0101" => d <= "11000110"; -- ##...##.
                when x"99" & "0110" => d <= "11000110"; -- ##...##.
                when x"99" & "0111" => d <= "11000110"; -- ##...##.
                when x"99" & "1000" => d <= "11000110"; -- ##...##.
                when x"99" & "1001" => d <= "11000110"; -- ##...##.
                when x"99" & "1010" => d <= "11000110"; -- ##...##.
                when x"99" & "1011" => d <= "01111100"; -- .#####..
                when x"99" & "1100" => d <= "00000000"; -- ........
                when x"99" & "1101" => d <= "00000000"; -- ........
                when x"99" & "1110" => d <= "00000000"; -- ........
                when x"99" & "1111" => d <= "00000000"; -- ........

                when x"9a" & "0000" => d <= "00000000"; -- ........
                when x"9a" & "0001" => d <= "11000110"; -- ##...##.
                when x"9a" & "0010" => d <= "00000000"; -- ........
                when x"9a" & "0011" => d <= "11000110"; -- ##...##.
                when x"9a" & "0100" => d <= "11000110"; -- ##...##.
                when x"9a" & "0101" => d <= "11000110"; -- ##...##.
                when x"9a" & "0110" => d <= "11000110"; -- ##...##.
                when x"9a" & "0111" => d <= "11000110"; -- ##...##.
                when x"9a" & "1000" => d <= "11000110"; -- ##...##.
                when x"9a" & "1001" => d <= "11000110"; -- ##...##.
                when x"9a" & "1010" => d <= "11000110"; -- ##...##.
                when x"9a" & "1011" => d <= "01111100"; -- .#####..
                when x"9a" & "1100" => d <= "00000000"; -- ........
                when x"9a" & "1101" => d <= "00000000"; -- ........
                when x"9a" & "1110" => d <= "00000000"; -- ........
                when x"9a" & "1111" => d <= "00000000"; -- ........

                when x"9b" & "0000" => d <= "00000000"; -- ........
                when x"9b" & "0001" => d <= "00011000"; -- ...##...
                when x"9b" & "0010" => d <= "00011000"; -- ...##...
                when x"9b" & "0011" => d <= "00111100"; -- ..####..
                when x"9b" & "0100" => d <= "01100110"; -- .##..##.
                when x"9b" & "0101" => d <= "01100000"; -- .##.....
                when x"9b" & "0110" => d <= "01100000"; -- .##.....
                when x"9b" & "0111" => d <= "01100000"; -- .##.....
                when x"9b" & "1000" => d <= "01100110"; -- .##..##.
                when x"9b" & "1001" => d <= "00111100"; -- ..####..
                when x"9b" & "1010" => d <= "00011000"; -- ...##...
                when x"9b" & "1011" => d <= "00011000"; -- ...##...
                when x"9b" & "1100" => d <= "00000000"; -- ........
                when x"9b" & "1101" => d <= "00000000"; -- ........
                when x"9b" & "1110" => d <= "00000000"; -- ........
                when x"9b" & "1111" => d <= "00000000"; -- ........

                when x"9c" & "0000" => d <= "00000000"; -- ........
                when x"9c" & "0001" => d <= "00111000"; -- ..###...
                when x"9c" & "0010" => d <= "01101100"; -- .##.##..
                when x"9c" & "0011" => d <= "01100100"; -- .##..#..
                when x"9c" & "0100" => d <= "01100000"; -- .##.....
                when x"9c" & "0101" => d <= "11110000"; -- ####....
                when x"9c" & "0110" => d <= "01100000"; -- .##.....
                when x"9c" & "0111" => d <= "01100000"; -- .##.....
                when x"9c" & "1000" => d <= "01100000"; -- .##.....
                when x"9c" & "1001" => d <= "01100000"; -- .##.....
                when x"9c" & "1010" => d <= "11100110"; -- ###..##.
                when x"9c" & "1011" => d <= "11111100"; -- ######..
                when x"9c" & "1100" => d <= "00000000"; -- ........
                when x"9c" & "1101" => d <= "00000000"; -- ........
                when x"9c" & "1110" => d <= "00000000"; -- ........
                when x"9c" & "1111" => d <= "00000000"; -- ........

                when x"9d" & "0000" => d <= "00000000"; -- ........
                when x"9d" & "0001" => d <= "00000000"; -- ........
                when x"9d" & "0010" => d <= "01100110"; -- .##..##.
                when x"9d" & "0011" => d <= "01100110"; -- .##..##.
                when x"9d" & "0100" => d <= "00111100"; -- ..####..
                when x"9d" & "0101" => d <= "00011000"; -- ...##...
                when x"9d" & "0110" => d <= "01111110"; -- .######.
                when x"9d" & "0111" => d <= "00011000"; -- ...##...
                when x"9d" & "1000" => d <= "01111110"; -- .######.
                when x"9d" & "1001" => d <= "00011000"; -- ...##...
                when x"9d" & "1010" => d <= "00011000"; -- ...##...
                when x"9d" & "1011" => d <= "00011000"; -- ...##...
                when x"9d" & "1100" => d <= "00000000"; -- ........
                when x"9d" & "1101" => d <= "00000000"; -- ........
                when x"9d" & "1110" => d <= "00000000"; -- ........
                when x"9d" & "1111" => d <= "00000000"; -- ........

                when x"9e" & "0000" => d <= "00000000"; -- ........
                when x"9e" & "0001" => d <= "11111000"; -- #####...
                when x"9e" & "0010" => d <= "11001100"; -- ##..##..
                when x"9e" & "0011" => d <= "11001100"; -- ##..##..
                when x"9e" & "0100" => d <= "11111000"; -- #####...
                when x"9e" & "0101" => d <= "11000100"; -- ##...#..
                when x"9e" & "0110" => d <= "11001100"; -- ##..##..
                when x"9e" & "0111" => d <= "11011110"; -- ##.####.
                when x"9e" & "1000" => d <= "11001100"; -- ##..##..
                when x"9e" & "1001" => d <= "11001100"; -- ##..##..
                when x"9e" & "1010" => d <= "11001100"; -- ##..##..
                when x"9e" & "1011" => d <= "11000110"; -- ##...##.
                when x"9e" & "1100" => d <= "00000000"; -- ........
                when x"9e" & "1101" => d <= "00000000"; -- ........
                when x"9e" & "1110" => d <= "00000000"; -- ........
                when x"9e" & "1111" => d <= "00000000"; -- ........

                when x"9f" & "0000" => d <= "00000000"; -- ........
                when x"9f" & "0001" => d <= "00001110"; -- ....###.
                when x"9f" & "0010" => d <= "00011011"; -- ...##.##
                when x"9f" & "0011" => d <= "00011000"; -- ...##...
                when x"9f" & "0100" => d <= "00011000"; -- ...##...
                when x"9f" & "0101" => d <= "00011000"; -- ...##...
                when x"9f" & "0110" => d <= "01111110"; -- .######.
                when x"9f" & "0111" => d <= "00011000"; -- ...##...
                when x"9f" & "1000" => d <= "00011000"; -- ...##...
                when x"9f" & "1001" => d <= "00011000"; -- ...##...
                when x"9f" & "1010" => d <= "00011000"; -- ...##...
                when x"9f" & "1011" => d <= "00011000"; -- ...##...
                when x"9f" & "1100" => d <= "11011000"; -- ##.##...
                when x"9f" & "1101" => d <= "01110000"; -- .###....
                when x"9f" & "1110" => d <= "00000000"; -- ........
                when x"9f" & "1111" => d <= "00000000"; -- ........

                when x"a0" & "0000" => d <= "00000000"; -- ........
                when x"a0" & "0001" => d <= "00011000"; -- ...##...
                when x"a0" & "0010" => d <= "00110000"; -- ..##....
                when x"a0" & "0011" => d <= "01100000"; -- .##.....
                when x"a0" & "0100" => d <= "00000000"; -- ........
                when x"a0" & "0101" => d <= "01111000"; -- .####...
                when x"a0" & "0110" => d <= "00001100"; -- ....##..
                when x"a0" & "0111" => d <= "01111100"; -- .#####..
                when x"a0" & "1000" => d <= "11001100"; -- ##..##..
                when x"a0" & "1001" => d <= "11001100"; -- ##..##..
                when x"a0" & "1010" => d <= "11001100"; -- ##..##..
                when x"a0" & "1011" => d <= "01110110"; -- .###.##.
                when x"a0" & "1100" => d <= "00000000"; -- ........
                when x"a0" & "1101" => d <= "00000000"; -- ........
                when x"a0" & "1110" => d <= "00000000"; -- ........
                when x"a0" & "1111" => d <= "00000000"; -- ........

                when x"a1" & "0000" => d <= "00000000"; -- ........
                when x"a1" & "0001" => d <= "00001100"; -- ....##..
                when x"a1" & "0010" => d <= "00011000"; -- ...##...
                when x"a1" & "0011" => d <= "00110000"; -- ..##....
                when x"a1" & "0100" => d <= "00000000"; -- ........
                when x"a1" & "0101" => d <= "00111000"; -- ..###...
                when x"a1" & "0110" => d <= "00011000"; -- ...##...
                when x"a1" & "0111" => d <= "00011000"; -- ...##...
                when x"a1" & "1000" => d <= "00011000"; -- ...##...
                when x"a1" & "1001" => d <= "00011000"; -- ...##...
                when x"a1" & "1010" => d <= "00011000"; -- ...##...
                when x"a1" & "1011" => d <= "00111100"; -- ..####..
                when x"a1" & "1100" => d <= "00000000"; -- ........
                when x"a1" & "1101" => d <= "00000000"; -- ........
                when x"a1" & "1110" => d <= "00000000"; -- ........
                when x"a1" & "1111" => d <= "00000000"; -- ........

                when x"a2" & "0000" => d <= "00000000"; -- ........
                when x"a2" & "0001" => d <= "00011000"; -- ...##...
                when x"a2" & "0010" => d <= "00110000"; -- ..##....
                when x"a2" & "0011" => d <= "01100000"; -- .##.....
                when x"a2" & "0100" => d <= "00000000"; -- ........
                when x"a2" & "0101" => d <= "01111100"; -- .#####..
                when x"a2" & "0110" => d <= "11000110"; -- ##...##.
                when x"a2" & "0111" => d <= "11000110"; -- ##...##.
                when x"a2" & "1000" => d <= "11000110"; -- ##...##.
                when x"a2" & "1001" => d <= "11000110"; -- ##...##.
                when x"a2" & "1010" => d <= "11000110"; -- ##...##.
                when x"a2" & "1011" => d <= "01111100"; -- .#####..
                when x"a2" & "1100" => d <= "00000000"; -- ........
                when x"a2" & "1101" => d <= "00000000"; -- ........
                when x"a2" & "1110" => d <= "00000000"; -- ........
                when x"a2" & "1111" => d <= "00000000"; -- ........

                when x"a3" & "0000" => d <= "00000000"; -- ........
                when x"a3" & "0001" => d <= "00011000"; -- ...##...
                when x"a3" & "0010" => d <= "00110000"; -- ..##....
                when x"a3" & "0011" => d <= "01100000"; -- .##.....
                when x"a3" & "0100" => d <= "00000000"; -- ........
                when x"a3" & "0101" => d <= "11001100"; -- ##..##..
                when x"a3" & "0110" => d <= "11001100"; -- ##..##..
                when x"a3" & "0111" => d <= "11001100"; -- ##..##..
                when x"a3" & "1000" => d <= "11001100"; -- ##..##..
                when x"a3" & "1001" => d <= "11001100"; -- ##..##..
                when x"a3" & "1010" => d <= "11001100"; -- ##..##..
                when x"a3" & "1011" => d <= "01110110"; -- .###.##.
                when x"a3" & "1100" => d <= "00000000"; -- ........
                when x"a3" & "1101" => d <= "00000000"; -- ........
                when x"a3" & "1110" => d <= "00000000"; -- ........
                when x"a3" & "1111" => d <= "00000000"; -- ........

                when x"a4" & "0000" => d <= "00000000"; -- ........
                when x"a4" & "0001" => d <= "00000000"; -- ........
                when x"a4" & "0010" => d <= "01110110"; -- .###.##.
                when x"a4" & "0011" => d <= "11011100"; -- ##.###..
                when x"a4" & "0100" => d <= "00000000"; -- ........
                when x"a4" & "0101" => d <= "11011100"; -- ##.###..
                when x"a4" & "0110" => d <= "01100110"; -- .##..##.
                when x"a4" & "0111" => d <= "01100110"; -- .##..##.
                when x"a4" & "1000" => d <= "01100110"; -- .##..##.
                when x"a4" & "1001" => d <= "01100110"; -- .##..##.
                when x"a4" & "1010" => d <= "01100110"; -- .##..##.
                when x"a4" & "1011" => d <= "01100110"; -- .##..##.
                when x"a4" & "1100" => d <= "00000000"; -- ........
                when x"a4" & "1101" => d <= "00000000"; -- ........
                when x"a4" & "1110" => d <= "00000000"; -- ........
                when x"a4" & "1111" => d <= "00000000"; -- ........

                when x"a5" & "0000" => d <= "01110110"; -- .###.##.
                when x"a5" & "0001" => d <= "11011100"; -- ##.###..
                when x"a5" & "0010" => d <= "00000000"; -- ........
                when x"a5" & "0011" => d <= "11000110"; -- ##...##.
                when x"a5" & "0100" => d <= "11100110"; -- ###..##.
                when x"a5" & "0101" => d <= "11110110"; -- ####.##.
                when x"a5" & "0110" => d <= "11111110"; -- #######.
                when x"a5" & "0111" => d <= "11011110"; -- ##.####.
                when x"a5" & "1000" => d <= "11001110"; -- ##..###.
                when x"a5" & "1001" => d <= "11000110"; -- ##...##.
                when x"a5" & "1010" => d <= "11000110"; -- ##...##.
                when x"a5" & "1011" => d <= "11000110"; -- ##...##.
                when x"a5" & "1100" => d <= "00000000"; -- ........
                when x"a5" & "1101" => d <= "00000000"; -- ........
                when x"a5" & "1110" => d <= "00000000"; -- ........
                when x"a5" & "1111" => d <= "00000000"; -- ........

                when x"a6" & "0000" => d <= "00000000"; -- ........
                when x"a6" & "0001" => d <= "00111100"; -- ..####..
                when x"a6" & "0010" => d <= "01101100"; -- .##.##..
                when x"a6" & "0011" => d <= "01101100"; -- .##.##..
                when x"a6" & "0100" => d <= "00111110"; -- ..#####.
                when x"a6" & "0101" => d <= "00000000"; -- ........
                when x"a6" & "0110" => d <= "01111110"; -- .######.
                when x"a6" & "0111" => d <= "00000000"; -- ........
                when x"a6" & "1000" => d <= "00000000"; -- ........
                when x"a6" & "1001" => d <= "00000000"; -- ........
                when x"a6" & "1010" => d <= "00000000"; -- ........
                when x"a6" & "1011" => d <= "00000000"; -- ........
                when x"a6" & "1100" => d <= "00000000"; -- ........
                when x"a6" & "1101" => d <= "00000000"; -- ........
                when x"a6" & "1110" => d <= "00000000"; -- ........
                when x"a6" & "1111" => d <= "00000000"; -- ........

                when x"a7" & "0000" => d <= "00000000"; -- ........
                when x"a7" & "0001" => d <= "00111000"; -- ..###...
                when x"a7" & "0010" => d <= "01101100"; -- .##.##..
                when x"a7" & "0011" => d <= "01101100"; -- .##.##..
                when x"a7" & "0100" => d <= "00111000"; -- ..###...
                when x"a7" & "0101" => d <= "00000000"; -- ........
                when x"a7" & "0110" => d <= "01111100"; -- .#####..
                when x"a7" & "0111" => d <= "00000000"; -- ........
                when x"a7" & "1000" => d <= "00000000"; -- ........
                when x"a7" & "1001" => d <= "00000000"; -- ........
                when x"a7" & "1010" => d <= "00000000"; -- ........
                when x"a7" & "1011" => d <= "00000000"; -- ........
                when x"a7" & "1100" => d <= "00000000"; -- ........
                when x"a7" & "1101" => d <= "00000000"; -- ........
                when x"a7" & "1110" => d <= "00000000"; -- ........
                when x"a7" & "1111" => d <= "00000000"; -- ........

                when x"a8" & "0000" => d <= "00000000"; -- ........
                when x"a8" & "0001" => d <= "00000000"; -- ........
                when x"a8" & "0010" => d <= "00110000"; -- ..##....
                when x"a8" & "0011" => d <= "00110000"; -- ..##....
                when x"a8" & "0100" => d <= "00000000"; -- ........
                when x"a8" & "0101" => d <= "00110000"; -- ..##....
                when x"a8" & "0110" => d <= "00110000"; -- ..##....
                when x"a8" & "0111" => d <= "01100000"; -- .##.....
                when x"a8" & "1000" => d <= "11000000"; -- ##......
                when x"a8" & "1001" => d <= "11000110"; -- ##...##.
                when x"a8" & "1010" => d <= "11000110"; -- ##...##.
                when x"a8" & "1011" => d <= "01111100"; -- .#####..
                when x"a8" & "1100" => d <= "00000000"; -- ........
                when x"a8" & "1101" => d <= "00000000"; -- ........
                when x"a8" & "1110" => d <= "00000000"; -- ........
                when x"a8" & "1111" => d <= "00000000"; -- ........

                when x"a9" & "0000" => d <= "00000000"; -- ........
                when x"a9" & "0001" => d <= "00000000"; -- ........
                when x"a9" & "0010" => d <= "00000000"; -- ........
                when x"a9" & "0011" => d <= "00000000"; -- ........
                when x"a9" & "0100" => d <= "00000000"; -- ........
                when x"a9" & "0101" => d <= "00000000"; -- ........
                when x"a9" & "0110" => d <= "11111110"; -- #######.
                when x"a9" & "0111" => d <= "11000000"; -- ##......
                when x"a9" & "1000" => d <= "11000000"; -- ##......
                when x"a9" & "1001" => d <= "11000000"; -- ##......
                when x"a9" & "1010" => d <= "11000000"; -- ##......
                when x"a9" & "1011" => d <= "00000000"; -- ........
                when x"a9" & "1100" => d <= "00000000"; -- ........
                when x"a9" & "1101" => d <= "00000000"; -- ........
                when x"a9" & "1110" => d <= "00000000"; -- ........
                when x"a9" & "1111" => d <= "00000000"; -- ........

                when x"aa" & "0000" => d <= "00000000"; -- ........
                when x"aa" & "0001" => d <= "00000000"; -- ........
                when x"aa" & "0010" => d <= "00000000"; -- ........
                when x"aa" & "0011" => d <= "00000000"; -- ........
                when x"aa" & "0100" => d <= "00000000"; -- ........
                when x"aa" & "0101" => d <= "00000000"; -- ........
                when x"aa" & "0110" => d <= "11111110"; -- #######.
                when x"aa" & "0111" => d <= "00000110"; -- .....##.
                when x"aa" & "1000" => d <= "00000110"; -- .....##.
                when x"aa" & "1001" => d <= "00000110"; -- .....##.
                when x"aa" & "1010" => d <= "00000110"; -- .....##.
                when x"aa" & "1011" => d <= "00000000"; -- ........
                when x"aa" & "1100" => d <= "00000000"; -- ........
                when x"aa" & "1101" => d <= "00000000"; -- ........
                when x"aa" & "1110" => d <= "00000000"; -- ........
                when x"aa" & "1111" => d <= "00000000"; -- ........

                when x"ab" & "0000" => d <= "00000000"; -- ........
                when x"ab" & "0001" => d <= "11000000"; -- ##......
                when x"ab" & "0010" => d <= "11000000"; -- ##......
                when x"ab" & "0011" => d <= "11000010"; -- ##....#.
                when x"ab" & "0100" => d <= "11000110"; -- ##...##.
                when x"ab" & "0101" => d <= "11001100"; -- ##..##..
                when x"ab" & "0110" => d <= "00011000"; -- ...##...
                when x"ab" & "0111" => d <= "00110000"; -- ..##....
                when x"ab" & "1000" => d <= "01100000"; -- .##.....
                when x"ab" & "1001" => d <= "11011100"; -- ##.###..
                when x"ab" & "1010" => d <= "10000110"; -- #....##.
                when x"ab" & "1011" => d <= "00001100"; -- ....##..
                when x"ab" & "1100" => d <= "00011000"; -- ...##...
                when x"ab" & "1101" => d <= "00111110"; -- ..#####.
                when x"ab" & "1110" => d <= "00000000"; -- ........
                when x"ab" & "1111" => d <= "00000000"; -- ........

                when x"ac" & "0000" => d <= "00000000"; -- ........
                when x"ac" & "0001" => d <= "11000000"; -- ##......
                when x"ac" & "0010" => d <= "11000000"; -- ##......
                when x"ac" & "0011" => d <= "11000010"; -- ##....#.
                when x"ac" & "0100" => d <= "11000110"; -- ##...##.
                when x"ac" & "0101" => d <= "11001100"; -- ##..##..
                when x"ac" & "0110" => d <= "00011000"; -- ...##...
                when x"ac" & "0111" => d <= "00110000"; -- ..##....
                when x"ac" & "1000" => d <= "01100110"; -- .##..##.
                when x"ac" & "1001" => d <= "11001110"; -- ##..###.
                when x"ac" & "1010" => d <= "10011110"; -- #..####.
                when x"ac" & "1011" => d <= "00111110"; -- ..#####.
                when x"ac" & "1100" => d <= "00000110"; -- .....##.
                when x"ac" & "1101" => d <= "00000110"; -- .....##.
                when x"ac" & "1110" => d <= "00000000"; -- ........
                when x"ac" & "1111" => d <= "00000000"; -- ........

                when x"ad" & "0000" => d <= "00000000"; -- ........
                when x"ad" & "0001" => d <= "00000000"; -- ........
                when x"ad" & "0010" => d <= "00011000"; -- ...##...
                when x"ad" & "0011" => d <= "00011000"; -- ...##...
                when x"ad" & "0100" => d <= "00000000"; -- ........
                when x"ad" & "0101" => d <= "00011000"; -- ...##...
                when x"ad" & "0110" => d <= "00011000"; -- ...##...
                when x"ad" & "0111" => d <= "00011000"; -- ...##...
                when x"ad" & "1000" => d <= "00111100"; -- ..####..
                when x"ad" & "1001" => d <= "00111100"; -- ..####..
                when x"ad" & "1010" => d <= "00111100"; -- ..####..
                when x"ad" & "1011" => d <= "00011000"; -- ...##...
                when x"ad" & "1100" => d <= "00000000"; -- ........
                when x"ad" & "1101" => d <= "00000000"; -- ........
                when x"ad" & "1110" => d <= "00000000"; -- ........
                when x"ad" & "1111" => d <= "00000000"; -- ........

                when x"ae" & "0000" => d <= "00000000"; -- ........
                when x"ae" & "0001" => d <= "00000000"; -- ........
                when x"ae" & "0010" => d <= "00000000"; -- ........
                when x"ae" & "0011" => d <= "00000000"; -- ........
                when x"ae" & "0100" => d <= "00000000"; -- ........
                when x"ae" & "0101" => d <= "00110110"; -- ..##.##.
                when x"ae" & "0110" => d <= "01101100"; -- .##.##..
                when x"ae" & "0111" => d <= "11011000"; -- ##.##...
                when x"ae" & "1000" => d <= "01101100"; -- .##.##..
                when x"ae" & "1001" => d <= "00110110"; -- ..##.##.
                when x"ae" & "1010" => d <= "00000000"; -- ........
                when x"ae" & "1011" => d <= "00000000"; -- ........
                when x"ae" & "1100" => d <= "00000000"; -- ........
                when x"ae" & "1101" => d <= "00000000"; -- ........
                when x"ae" & "1110" => d <= "00000000"; -- ........
                when x"ae" & "1111" => d <= "00000000"; -- ........

                when x"af" & "0000" => d <= "00000000"; -- ........
                when x"af" & "0001" => d <= "00000000"; -- ........
                when x"af" & "0010" => d <= "00000000"; -- ........
                when x"af" & "0011" => d <= "00000000"; -- ........
                when x"af" & "0100" => d <= "00000000"; -- ........
                when x"af" & "0101" => d <= "11011000"; -- ##.##...
                when x"af" & "0110" => d <= "01101100"; -- .##.##..
                when x"af" & "0111" => d <= "00110110"; -- ..##.##.
                when x"af" & "1000" => d <= "01101100"; -- .##.##..
                when x"af" & "1001" => d <= "11011000"; -- ##.##...
                when x"af" & "1010" => d <= "00000000"; -- ........
                when x"af" & "1011" => d <= "00000000"; -- ........
                when x"af" & "1100" => d <= "00000000"; -- ........
                when x"af" & "1101" => d <= "00000000"; -- ........
                when x"af" & "1110" => d <= "00000000"; -- ........
                when x"af" & "1111" => d <= "00000000"; -- ........

                when x"b0" & "0000" => d <= "00010001"; -- ...#...#
                when x"b0" & "0001" => d <= "01000100"; -- .#...#..
                when x"b0" & "0010" => d <= "00010001"; -- ...#...#
                when x"b0" & "0011" => d <= "01000100"; -- .#...#..
                when x"b0" & "0100" => d <= "00010001"; -- ...#...#
                when x"b0" & "0101" => d <= "01000100"; -- .#...#..
                when x"b0" & "0110" => d <= "00010001"; -- ...#...#
                when x"b0" & "0111" => d <= "01000100"; -- .#...#..
                when x"b0" & "1000" => d <= "00010001"; -- ...#...#
                when x"b0" & "1001" => d <= "01000100"; -- .#...#..
                when x"b0" & "1010" => d <= "00010001"; -- ...#...#
                when x"b0" & "1011" => d <= "01000100"; -- .#...#..
                when x"b0" & "1100" => d <= "00010001"; -- ...#...#
                when x"b0" & "1101" => d <= "01000100"; -- .#...#..
                when x"b0" & "1110" => d <= "00010001"; -- ...#...#
                when x"b0" & "1111" => d <= "01000100"; -- .#...#..

                when x"b1" & "0000" => d <= "01010101"; -- .#.#.#.#
                when x"b1" & "0001" => d <= "10101010"; -- #.#.#.#.
                when x"b1" & "0010" => d <= "01010101"; -- .#.#.#.#
                when x"b1" & "0011" => d <= "10101010"; -- #.#.#.#.
                when x"b1" & "0100" => d <= "01010101"; -- .#.#.#.#
                when x"b1" & "0101" => d <= "10101010"; -- #.#.#.#.
                when x"b1" & "0110" => d <= "01010101"; -- .#.#.#.#
                when x"b1" & "0111" => d <= "10101010"; -- #.#.#.#.
                when x"b1" & "1000" => d <= "01010101"; -- .#.#.#.#
                when x"b1" & "1001" => d <= "10101010"; -- #.#.#.#.
                when x"b1" & "1010" => d <= "01010101"; -- .#.#.#.#
                when x"b1" & "1011" => d <= "10101010"; -- #.#.#.#.
                when x"b1" & "1100" => d <= "01010101"; -- .#.#.#.#
                when x"b1" & "1101" => d <= "10101010"; -- #.#.#.#.
                when x"b1" & "1110" => d <= "01010101"; -- .#.#.#.#
                when x"b1" & "1111" => d <= "10101010"; -- #.#.#.#.

                when x"b2" & "0000" => d <= "11011101"; -- ##.###.#
                when x"b2" & "0001" => d <= "01110111"; -- .###.###
                when x"b2" & "0010" => d <= "11011101"; -- ##.###.#
                when x"b2" & "0011" => d <= "01110111"; -- .###.###
                when x"b2" & "0100" => d <= "11011101"; -- ##.###.#
                when x"b2" & "0101" => d <= "01110111"; -- .###.###
                when x"b2" & "0110" => d <= "11011101"; -- ##.###.#
                when x"b2" & "0111" => d <= "01110111"; -- .###.###
                when x"b2" & "1000" => d <= "11011101"; -- ##.###.#
                when x"b2" & "1001" => d <= "01110111"; -- .###.###
                when x"b2" & "1010" => d <= "11011101"; -- ##.###.#
                when x"b2" & "1011" => d <= "01110111"; -- .###.###
                when x"b2" & "1100" => d <= "11011101"; -- ##.###.#
                when x"b2" & "1101" => d <= "01110111"; -- .###.###
                when x"b2" & "1110" => d <= "11011101"; -- ##.###.#
                when x"b2" & "1111" => d <= "01110111"; -- .###.###

                when x"b3" & "0000" => d <= "00011000"; -- ...##...
                when x"b3" & "0001" => d <= "00011000"; -- ...##...
                when x"b3" & "0010" => d <= "00011000"; -- ...##...
                when x"b3" & "0011" => d <= "00011000"; -- ...##...
                when x"b3" & "0100" => d <= "00011000"; -- ...##...
                when x"b3" & "0101" => d <= "00011000"; -- ...##...
                when x"b3" & "0110" => d <= "00011000"; -- ...##...
                when x"b3" & "0111" => d <= "00011000"; -- ...##...
                when x"b3" & "1000" => d <= "00011000"; -- ...##...
                when x"b3" & "1001" => d <= "00011000"; -- ...##...
                when x"b3" & "1010" => d <= "00011000"; -- ...##...
                when x"b3" & "1011" => d <= "00011000"; -- ...##...
                when x"b3" & "1100" => d <= "00011000"; -- ...##...
                when x"b3" & "1101" => d <= "00011000"; -- ...##...
                when x"b3" & "1110" => d <= "00011000"; -- ...##...
                when x"b3" & "1111" => d <= "00011000"; -- ...##...

                when x"b4" & "0000" => d <= "00011000"; -- ...##...
                when x"b4" & "0001" => d <= "00011000"; -- ...##...
                when x"b4" & "0010" => d <= "00011000"; -- ...##...
                when x"b4" & "0011" => d <= "00011000"; -- ...##...
                when x"b4" & "0100" => d <= "00011000"; -- ...##...
                when x"b4" & "0101" => d <= "00011000"; -- ...##...
                when x"b4" & "0110" => d <= "00011000"; -- ...##...
                when x"b4" & "0111" => d <= "11111000"; -- #####...
                when x"b4" & "1000" => d <= "00011000"; -- ...##...
                when x"b4" & "1001" => d <= "00011000"; -- ...##...
                when x"b4" & "1010" => d <= "00011000"; -- ...##...
                when x"b4" & "1011" => d <= "00011000"; -- ...##...
                when x"b4" & "1100" => d <= "00011000"; -- ...##...
                when x"b4" & "1101" => d <= "00011000"; -- ...##...
                when x"b4" & "1110" => d <= "00011000"; -- ...##...
                when x"b4" & "1111" => d <= "00011000"; -- ...##...

                when x"b5" & "0000" => d <= "00011000"; -- ...##...
                when x"b5" & "0001" => d <= "00011000"; -- ...##...
                when x"b5" & "0010" => d <= "00011000"; -- ...##...
                when x"b5" & "0011" => d <= "00011000"; -- ...##...
                when x"b5" & "0100" => d <= "00011000"; -- ...##...
                when x"b5" & "0101" => d <= "11111000"; -- #####...
                when x"b5" & "0110" => d <= "00011000"; -- ...##...
                when x"b5" & "0111" => d <= "11111000"; -- #####...
                when x"b5" & "1000" => d <= "00011000"; -- ...##...
                when x"b5" & "1001" => d <= "00011000"; -- ...##...
                when x"b5" & "1010" => d <= "00011000"; -- ...##...
                when x"b5" & "1011" => d <= "00011000"; -- ...##...
                when x"b5" & "1100" => d <= "00011000"; -- ...##...
                when x"b5" & "1101" => d <= "00011000"; -- ...##...
                when x"b5" & "1110" => d <= "00011000"; -- ...##...
                when x"b5" & "1111" => d <= "00011000"; -- ...##...

                when x"b6" & "0000" => d <= "00110110"; -- ..##.##.
                when x"b6" & "0001" => d <= "00110110"; -- ..##.##.
                when x"b6" & "0010" => d <= "00110110"; -- ..##.##.
                when x"b6" & "0011" => d <= "00110110"; -- ..##.##.
                when x"b6" & "0100" => d <= "00110110"; -- ..##.##.
                when x"b6" & "0101" => d <= "00110110"; -- ..##.##.
                when x"b6" & "0110" => d <= "00110110"; -- ..##.##.
                when x"b6" & "0111" => d <= "11110110"; -- ####.##.
                when x"b6" & "1000" => d <= "00110110"; -- ..##.##.
                when x"b6" & "1001" => d <= "00110110"; -- ..##.##.
                when x"b6" & "1010" => d <= "00110110"; -- ..##.##.
                when x"b6" & "1011" => d <= "00110110"; -- ..##.##.
                when x"b6" & "1100" => d <= "00110110"; -- ..##.##.
                when x"b6" & "1101" => d <= "00110110"; -- ..##.##.
                when x"b6" & "1110" => d <= "00110110"; -- ..##.##.
                when x"b6" & "1111" => d <= "00110110"; -- ..##.##.

                when x"b7" & "0000" => d <= "00000000"; -- ........
                when x"b7" & "0001" => d <= "00000000"; -- ........
                when x"b7" & "0010" => d <= "00000000"; -- ........
                when x"b7" & "0011" => d <= "00000000"; -- ........
                when x"b7" & "0100" => d <= "00000000"; -- ........
                when x"b7" & "0101" => d <= "00000000"; -- ........
                when x"b7" & "0110" => d <= "00000000"; -- ........
                when x"b7" & "0111" => d <= "11111110"; -- #######.
                when x"b7" & "1000" => d <= "00110110"; -- ..##.##.
                when x"b7" & "1001" => d <= "00110110"; -- ..##.##.
                when x"b7" & "1010" => d <= "00110110"; -- ..##.##.
                when x"b7" & "1011" => d <= "00110110"; -- ..##.##.
                when x"b7" & "1100" => d <= "00110110"; -- ..##.##.
                when x"b7" & "1101" => d <= "00110110"; -- ..##.##.
                when x"b7" & "1110" => d <= "00110110"; -- ..##.##.
                when x"b7" & "1111" => d <= "00110110"; -- ..##.##.

                when x"b8" & "0000" => d <= "00000000"; -- ........
                when x"b8" & "0001" => d <= "00000000"; -- ........
                when x"b8" & "0010" => d <= "00000000"; -- ........
                when x"b8" & "0011" => d <= "00000000"; -- ........
                when x"b8" & "0100" => d <= "00000000"; -- ........
                when x"b8" & "0101" => d <= "11111000"; -- #####...
                when x"b8" & "0110" => d <= "00011000"; -- ...##...
                when x"b8" & "0111" => d <= "11111000"; -- #####...
                when x"b8" & "1000" => d <= "00011000"; -- ...##...
                when x"b8" & "1001" => d <= "00011000"; -- ...##...
                when x"b8" & "1010" => d <= "00011000"; -- ...##...
                when x"b8" & "1011" => d <= "00011000"; -- ...##...
                when x"b8" & "1100" => d <= "00011000"; -- ...##...
                when x"b8" & "1101" => d <= "00011000"; -- ...##...
                when x"b8" & "1110" => d <= "00011000"; -- ...##...
                when x"b8" & "1111" => d <= "00011000"; -- ...##...

                when x"b9" & "0000" => d <= "00110110"; -- ..##.##.
                when x"b9" & "0001" => d <= "00110110"; -- ..##.##.
                when x"b9" & "0010" => d <= "00110110"; -- ..##.##.
                when x"b9" & "0011" => d <= "00110110"; -- ..##.##.
                when x"b9" & "0100" => d <= "00110110"; -- ..##.##.
                when x"b9" & "0101" => d <= "11110110"; -- ####.##.
                when x"b9" & "0110" => d <= "00000110"; -- .....##.
                when x"b9" & "0111" => d <= "11110110"; -- ####.##.
                when x"b9" & "1000" => d <= "00110110"; -- ..##.##.
                when x"b9" & "1001" => d <= "00110110"; -- ..##.##.
                when x"b9" & "1010" => d <= "00110110"; -- ..##.##.
                when x"b9" & "1011" => d <= "00110110"; -- ..##.##.
                when x"b9" & "1100" => d <= "00110110"; -- ..##.##.
                when x"b9" & "1101" => d <= "00110110"; -- ..##.##.
                when x"b9" & "1110" => d <= "00110110"; -- ..##.##.
                when x"b9" & "1111" => d <= "00110110"; -- ..##.##.

                when x"ba" & "0000" => d <= "00110110"; -- ..##.##.
                when x"ba" & "0001" => d <= "00110110"; -- ..##.##.
                when x"ba" & "0010" => d <= "00110110"; -- ..##.##.
                when x"ba" & "0011" => d <= "00110110"; -- ..##.##.
                when x"ba" & "0100" => d <= "00110110"; -- ..##.##.
                when x"ba" & "0101" => d <= "00110110"; -- ..##.##.
                when x"ba" & "0110" => d <= "00110110"; -- ..##.##.
                when x"ba" & "0111" => d <= "00110110"; -- ..##.##.
                when x"ba" & "1000" => d <= "00110110"; -- ..##.##.
                when x"ba" & "1001" => d <= "00110110"; -- ..##.##.
                when x"ba" & "1010" => d <= "00110110"; -- ..##.##.
                when x"ba" & "1011" => d <= "00110110"; -- ..##.##.
                when x"ba" & "1100" => d <= "00110110"; -- ..##.##.
                when x"ba" & "1101" => d <= "00110110"; -- ..##.##.
                when x"ba" & "1110" => d <= "00110110"; -- ..##.##.
                when x"ba" & "1111" => d <= "00110110"; -- ..##.##.

                when x"bb" & "0000" => d <= "00000000"; -- ........
                when x"bb" & "0001" => d <= "00000000"; -- ........
                when x"bb" & "0010" => d <= "00000000"; -- ........
                when x"bb" & "0011" => d <= "00000000"; -- ........
                when x"bb" & "0100" => d <= "00000000"; -- ........
                when x"bb" & "0101" => d <= "11111110"; -- #######.
                when x"bb" & "0110" => d <= "00000110"; -- .....##.
                when x"bb" & "0111" => d <= "11110110"; -- ####.##.
                when x"bb" & "1000" => d <= "00110110"; -- ..##.##.
                when x"bb" & "1001" => d <= "00110110"; -- ..##.##.
                when x"bb" & "1010" => d <= "00110110"; -- ..##.##.
                when x"bb" & "1011" => d <= "00110110"; -- ..##.##.
                when x"bb" & "1100" => d <= "00110110"; -- ..##.##.
                when x"bb" & "1101" => d <= "00110110"; -- ..##.##.
                when x"bb" & "1110" => d <= "00110110"; -- ..##.##.
                when x"bb" & "1111" => d <= "00110110"; -- ..##.##.

                when x"bc" & "0000" => d <= "00110110"; -- ..##.##.
                when x"bc" & "0001" => d <= "00110110"; -- ..##.##.
                when x"bc" & "0010" => d <= "00110110"; -- ..##.##.
                when x"bc" & "0011" => d <= "00110110"; -- ..##.##.
                when x"bc" & "0100" => d <= "00110110"; -- ..##.##.
                when x"bc" & "0101" => d <= "11110110"; -- ####.##.
                when x"bc" & "0110" => d <= "00000110"; -- .....##.
                when x"bc" & "0111" => d <= "11111110"; -- #######.
                when x"bc" & "1000" => d <= "00000000"; -- ........
                when x"bc" & "1001" => d <= "00000000"; -- ........
                when x"bc" & "1010" => d <= "00000000"; -- ........
                when x"bc" & "1011" => d <= "00000000"; -- ........
                when x"bc" & "1100" => d <= "00000000"; -- ........
                when x"bc" & "1101" => d <= "00000000"; -- ........
                when x"bc" & "1110" => d <= "00000000"; -- ........
                when x"bc" & "1111" => d <= "00000000"; -- ........

                when x"bd" & "0000" => d <= "00110110"; -- ..##.##.
                when x"bd" & "0001" => d <= "00110110"; -- ..##.##.
                when x"bd" & "0010" => d <= "00110110"; -- ..##.##.
                when x"bd" & "0011" => d <= "00110110"; -- ..##.##.
                when x"bd" & "0100" => d <= "00110110"; -- ..##.##.
                when x"bd" & "0101" => d <= "00110110"; -- ..##.##.
                when x"bd" & "0110" => d <= "00110110"; -- ..##.##.
                when x"bd" & "0111" => d <= "11111110"; -- #######.
                when x"bd" & "1000" => d <= "00000000"; -- ........
                when x"bd" & "1001" => d <= "00000000"; -- ........
                when x"bd" & "1010" => d <= "00000000"; -- ........
                when x"bd" & "1011" => d <= "00000000"; -- ........
                when x"bd" & "1100" => d <= "00000000"; -- ........
                when x"bd" & "1101" => d <= "00000000"; -- ........
                when x"bd" & "1110" => d <= "00000000"; -- ........
                when x"bd" & "1111" => d <= "00000000"; -- ........

                when x"be" & "0000" => d <= "00011000"; -- ...##...
                when x"be" & "0001" => d <= "00011000"; -- ...##...
                when x"be" & "0010" => d <= "00011000"; -- ...##...
                when x"be" & "0011" => d <= "00011000"; -- ...##...
                when x"be" & "0100" => d <= "00011000"; -- ...##...
                when x"be" & "0101" => d <= "11111000"; -- #####...
                when x"be" & "0110" => d <= "00011000"; -- ...##...
                when x"be" & "0111" => d <= "11111000"; -- #####...
                when x"be" & "1000" => d <= "00000000"; -- ........
                when x"be" & "1001" => d <= "00000000"; -- ........
                when x"be" & "1010" => d <= "00000000"; -- ........
                when x"be" & "1011" => d <= "00000000"; -- ........
                when x"be" & "1100" => d <= "00000000"; -- ........
                when x"be" & "1101" => d <= "00000000"; -- ........
                when x"be" & "1110" => d <= "00000000"; -- ........
                when x"be" & "1111" => d <= "00000000"; -- ........

                when x"bf" & "0000" => d <= "00000000"; -- ........
                when x"bf" & "0001" => d <= "00000000"; -- ........
                when x"bf" & "0010" => d <= "00000000"; -- ........
                when x"bf" & "0011" => d <= "00000000"; -- ........
                when x"bf" & "0100" => d <= "00000000"; -- ........
                when x"bf" & "0101" => d <= "00000000"; -- ........
                when x"bf" & "0110" => d <= "00000000"; -- ........
                when x"bf" & "0111" => d <= "11111000"; -- #####...
                when x"bf" & "1000" => d <= "00011000"; -- ...##...
                when x"bf" & "1001" => d <= "00011000"; -- ...##...
                when x"bf" & "1010" => d <= "00011000"; -- ...##...
                when x"bf" & "1011" => d <= "00011000"; -- ...##...
                when x"bf" & "1100" => d <= "00011000"; -- ...##...
                when x"bf" & "1101" => d <= "00011000"; -- ...##...
                when x"bf" & "1110" => d <= "00011000"; -- ...##...
                when x"bf" & "1111" => d <= "00011000"; -- ...##...

                when x"c0" & "0000" => d <= "00011000"; -- ...##...
                when x"c0" & "0001" => d <= "00011000"; -- ...##...
                when x"c0" & "0010" => d <= "00011000"; -- ...##...
                when x"c0" & "0011" => d <= "00011000"; -- ...##...
                when x"c0" & "0100" => d <= "00011000"; -- ...##...
                when x"c0" & "0101" => d <= "00011000"; -- ...##...
                when x"c0" & "0110" => d <= "00011000"; -- ...##...
                when x"c0" & "0111" => d <= "00011111"; -- ...#####
                when x"c0" & "1000" => d <= "00000000"; -- ........
                when x"c0" & "1001" => d <= "00000000"; -- ........
                when x"c0" & "1010" => d <= "00000000"; -- ........
                when x"c0" & "1011" => d <= "00000000"; -- ........
                when x"c0" & "1100" => d <= "00000000"; -- ........
                when x"c0" & "1101" => d <= "00000000"; -- ........
                when x"c0" & "1110" => d <= "00000000"; -- ........
                when x"c0" & "1111" => d <= "00000000"; -- ........

                when x"c1" & "0000" => d <= "00011000"; -- ...##...
                when x"c1" & "0001" => d <= "00011000"; -- ...##...
                when x"c1" & "0010" => d <= "00011000"; -- ...##...
                when x"c1" & "0011" => d <= "00011000"; -- ...##...
                when x"c1" & "0100" => d <= "00011000"; -- ...##...
                when x"c1" & "0101" => d <= "00011000"; -- ...##...
                when x"c1" & "0110" => d <= "00011000"; -- ...##...
                when x"c1" & "0111" => d <= "11111111"; -- ########
                when x"c1" & "1000" => d <= "00000000"; -- ........
                when x"c1" & "1001" => d <= "00000000"; -- ........
                when x"c1" & "1010" => d <= "00000000"; -- ........
                when x"c1" & "1011" => d <= "00000000"; -- ........
                when x"c1" & "1100" => d <= "00000000"; -- ........
                when x"c1" & "1101" => d <= "00000000"; -- ........
                when x"c1" & "1110" => d <= "00000000"; -- ........
                when x"c1" & "1111" => d <= "00000000"; -- ........

                when x"c2" & "0000" => d <= "00000000"; -- ........
                when x"c2" & "0001" => d <= "00000000"; -- ........
                when x"c2" & "0010" => d <= "00000000"; -- ........
                when x"c2" & "0011" => d <= "00000000"; -- ........
                when x"c2" & "0100" => d <= "00000000"; -- ........
                when x"c2" & "0101" => d <= "00000000"; -- ........
                when x"c2" & "0110" => d <= "00000000"; -- ........
                when x"c2" & "0111" => d <= "11111111"; -- ########
                when x"c2" & "1000" => d <= "00011000"; -- ...##...
                when x"c2" & "1001" => d <= "00011000"; -- ...##...
                when x"c2" & "1010" => d <= "00011000"; -- ...##...
                when x"c2" & "1011" => d <= "00011000"; -- ...##...
                when x"c2" & "1100" => d <= "00011000"; -- ...##...
                when x"c2" & "1101" => d <= "00011000"; -- ...##...
                when x"c2" & "1110" => d <= "00011000"; -- ...##...
                when x"c2" & "1111" => d <= "00011000"; -- ...##...

                when x"c3" & "0000" => d <= "00011000"; -- ...##...
                when x"c3" & "0001" => d <= "00011000"; -- ...##...
                when x"c3" & "0010" => d <= "00011000"; -- ...##...
                when x"c3" & "0011" => d <= "00011000"; -- ...##...
                when x"c3" & "0100" => d <= "00011000"; -- ...##...
                when x"c3" & "0101" => d <= "00011000"; -- ...##...
                when x"c3" & "0110" => d <= "00011000"; -- ...##...
                when x"c3" & "0111" => d <= "00011111"; -- ...#####
                when x"c3" & "1000" => d <= "00011000"; -- ...##...
                when x"c3" & "1001" => d <= "00011000"; -- ...##...
                when x"c3" & "1010" => d <= "00011000"; -- ...##...
                when x"c3" & "1011" => d <= "00011000"; -- ...##...
                when x"c3" & "1100" => d <= "00011000"; -- ...##...
                when x"c3" & "1101" => d <= "00011000"; -- ...##...
                when x"c3" & "1110" => d <= "00011000"; -- ...##...
                when x"c3" & "1111" => d <= "00011000"; -- ...##...

                when x"c4" & "0000" => d <= "00000000"; -- ........
                when x"c4" & "0001" => d <= "00000000"; -- ........
                when x"c4" & "0010" => d <= "00000000"; -- ........
                when x"c4" & "0011" => d <= "00000000"; -- ........
                when x"c4" & "0100" => d <= "00000000"; -- ........
                when x"c4" & "0101" => d <= "00000000"; -- ........
                when x"c4" & "0110" => d <= "00000000"; -- ........
                when x"c4" & "0111" => d <= "11111111"; -- ########
                when x"c4" & "1000" => d <= "00000000"; -- ........
                when x"c4" & "1001" => d <= "00000000"; -- ........
                when x"c4" & "1010" => d <= "00000000"; -- ........
                when x"c4" & "1011" => d <= "00000000"; -- ........
                when x"c4" & "1100" => d <= "00000000"; -- ........
                when x"c4" & "1101" => d <= "00000000"; -- ........
                when x"c4" & "1110" => d <= "00000000"; -- ........
                when x"c4" & "1111" => d <= "00000000"; -- ........

                when x"c5" & "0000" => d <= "00011000"; -- ...##...
                when x"c5" & "0001" => d <= "00011000"; -- ...##...
                when x"c5" & "0010" => d <= "00011000"; -- ...##...
                when x"c5" & "0011" => d <= "00011000"; -- ...##...
                when x"c5" & "0100" => d <= "00011000"; -- ...##...
                when x"c5" & "0101" => d <= "00011000"; -- ...##...
                when x"c5" & "0110" => d <= "00011000"; -- ...##...
                when x"c5" & "0111" => d <= "11111111"; -- ########
                when x"c5" & "1000" => d <= "00011000"; -- ...##...
                when x"c5" & "1001" => d <= "00011000"; -- ...##...
                when x"c5" & "1010" => d <= "00011000"; -- ...##...
                when x"c5" & "1011" => d <= "00011000"; -- ...##...
                when x"c5" & "1100" => d <= "00011000"; -- ...##...
                when x"c5" & "1101" => d <= "00011000"; -- ...##...
                when x"c5" & "1110" => d <= "00011000"; -- ...##...
                when x"c5" & "1111" => d <= "00011000"; -- ...##...

                when x"c6" & "0000" => d <= "00011000"; -- ...##...
                when x"c6" & "0001" => d <= "00011000"; -- ...##...
                when x"c6" & "0010" => d <= "00011000"; -- ...##...
                when x"c6" & "0011" => d <= "00011000"; -- ...##...
                when x"c6" & "0100" => d <= "00011000"; -- ...##...
                when x"c6" & "0101" => d <= "00011111"; -- ...#####
                when x"c6" & "0110" => d <= "00011000"; -- ...##...
                when x"c6" & "0111" => d <= "00011111"; -- ...#####
                when x"c6" & "1000" => d <= "00011000"; -- ...##...
                when x"c6" & "1001" => d <= "00011000"; -- ...##...
                when x"c6" & "1010" => d <= "00011000"; -- ...##...
                when x"c6" & "1011" => d <= "00011000"; -- ...##...
                when x"c6" & "1100" => d <= "00011000"; -- ...##...
                when x"c6" & "1101" => d <= "00011000"; -- ...##...
                when x"c6" & "1110" => d <= "00011000"; -- ...##...
                when x"c6" & "1111" => d <= "00011000"; -- ...##...

                when x"c7" & "0000" => d <= "00110110"; -- ..##.##.
                when x"c7" & "0001" => d <= "00110110"; -- ..##.##.
                when x"c7" & "0010" => d <= "00110110"; -- ..##.##.
                when x"c7" & "0011" => d <= "00110110"; -- ..##.##.
                when x"c7" & "0100" => d <= "00110110"; -- ..##.##.
                when x"c7" & "0101" => d <= "00110110"; -- ..##.##.
                when x"c7" & "0110" => d <= "00110110"; -- ..##.##.
                when x"c7" & "0111" => d <= "00110111"; -- ..##.###
                when x"c7" & "1000" => d <= "00110110"; -- ..##.##.
                when x"c7" & "1001" => d <= "00110110"; -- ..##.##.
                when x"c7" & "1010" => d <= "00110110"; -- ..##.##.
                when x"c7" & "1011" => d <= "00110110"; -- ..##.##.
                when x"c7" & "1100" => d <= "00110110"; -- ..##.##.
                when x"c7" & "1101" => d <= "00110110"; -- ..##.##.
                when x"c7" & "1110" => d <= "00110110"; -- ..##.##.
                when x"c7" & "1111" => d <= "00110110"; -- ..##.##.

                when x"c8" & "0000" => d <= "00110110"; -- ..##.##.
                when x"c8" & "0001" => d <= "00110110"; -- ..##.##.
                when x"c8" & "0010" => d <= "00110110"; -- ..##.##.
                when x"c8" & "0011" => d <= "00110110"; -- ..##.##.
                when x"c8" & "0100" => d <= "00110110"; -- ..##.##.
                when x"c8" & "0101" => d <= "00110111"; -- ..##.###
                when x"c8" & "0110" => d <= "00110000"; -- ..##....
                when x"c8" & "0111" => d <= "00111111"; -- ..######
                when x"c8" & "1000" => d <= "00000000"; -- ........
                when x"c8" & "1001" => d <= "00000000"; -- ........
                when x"c8" & "1010" => d <= "00000000"; -- ........
                when x"c8" & "1011" => d <= "00000000"; -- ........
                when x"c8" & "1100" => d <= "00000000"; -- ........
                when x"c8" & "1101" => d <= "00000000"; -- ........
                when x"c8" & "1110" => d <= "00000000"; -- ........
                when x"c8" & "1111" => d <= "00000000"; -- ........

                when x"c9" & "0000" => d <= "00000000"; -- ........
                when x"c9" & "0001" => d <= "00000000"; -- ........
                when x"c9" & "0010" => d <= "00000000"; -- ........
                when x"c9" & "0011" => d <= "00000000"; -- ........
                when x"c9" & "0100" => d <= "00000000"; -- ........
                when x"c9" & "0101" => d <= "00111111"; -- ..######
                when x"c9" & "0110" => d <= "00110000"; -- ..##....
                when x"c9" & "0111" => d <= "00110111"; -- ..##.###
                when x"c9" & "1000" => d <= "00110110"; -- ..##.##.
                when x"c9" & "1001" => d <= "00110110"; -- ..##.##.
                when x"c9" & "1010" => d <= "00110110"; -- ..##.##.
                when x"c9" & "1011" => d <= "00110110"; -- ..##.##.
                when x"c9" & "1100" => d <= "00110110"; -- ..##.##.
                when x"c9" & "1101" => d <= "00110110"; -- ..##.##.
                when x"c9" & "1110" => d <= "00110110"; -- ..##.##.
                when x"c9" & "1111" => d <= "00110110"; -- ..##.##.

                when x"ca" & "0000" => d <= "00110110"; -- ..##.##.
                when x"ca" & "0001" => d <= "00110110"; -- ..##.##.
                when x"ca" & "0010" => d <= "00110110"; -- ..##.##.
                when x"ca" & "0011" => d <= "00110110"; -- ..##.##.
                when x"ca" & "0100" => d <= "00110110"; -- ..##.##.
                when x"ca" & "0101" => d <= "11110111"; -- ####.###
                when x"ca" & "0110" => d <= "00000000"; -- ........
                when x"ca" & "0111" => d <= "11111111"; -- ########
                when x"ca" & "1000" => d <= "00000000"; -- ........
                when x"ca" & "1001" => d <= "00000000"; -- ........
                when x"ca" & "1010" => d <= "00000000"; -- ........
                when x"ca" & "1011" => d <= "00000000"; -- ........
                when x"ca" & "1100" => d <= "00000000"; -- ........
                when x"ca" & "1101" => d <= "00000000"; -- ........
                when x"ca" & "1110" => d <= "00000000"; -- ........
                when x"ca" & "1111" => d <= "00000000"; -- ........

                when x"cb" & "0000" => d <= "00000000"; -- ........
                when x"cb" & "0001" => d <= "00000000"; -- ........
                when x"cb" & "0010" => d <= "00000000"; -- ........
                when x"cb" & "0011" => d <= "00000000"; -- ........
                when x"cb" & "0100" => d <= "00000000"; -- ........
                when x"cb" & "0101" => d <= "11111111"; -- ########
                when x"cb" & "0110" => d <= "00000000"; -- ........
                when x"cb" & "0111" => d <= "11110111"; -- ####.###
                when x"cb" & "1000" => d <= "00110110"; -- ..##.##.
                when x"cb" & "1001" => d <= "00110110"; -- ..##.##.
                when x"cb" & "1010" => d <= "00110110"; -- ..##.##.
                when x"cb" & "1011" => d <= "00110110"; -- ..##.##.
                when x"cb" & "1100" => d <= "00110110"; -- ..##.##.
                when x"cb" & "1101" => d <= "00110110"; -- ..##.##.
                when x"cb" & "1110" => d <= "00110110"; -- ..##.##.
                when x"cb" & "1111" => d <= "00110110"; -- ..##.##.

                when x"cc" & "0000" => d <= "00110110"; -- ..##.##.
                when x"cc" & "0001" => d <= "00110110"; -- ..##.##.
                when x"cc" & "0010" => d <= "00110110"; -- ..##.##.
                when x"cc" & "0011" => d <= "00110110"; -- ..##.##.
                when x"cc" & "0100" => d <= "00110110"; -- ..##.##.
                when x"cc" & "0101" => d <= "00110111"; -- ..##.###
                when x"cc" & "0110" => d <= "00110000"; -- ..##....
                when x"cc" & "0111" => d <= "00110111"; -- ..##.###
                when x"cc" & "1000" => d <= "00110110"; -- ..##.##.
                when x"cc" & "1001" => d <= "00110110"; -- ..##.##.
                when x"cc" & "1010" => d <= "00110110"; -- ..##.##.
                when x"cc" & "1011" => d <= "00110110"; -- ..##.##.
                when x"cc" & "1100" => d <= "00110110"; -- ..##.##.
                when x"cc" & "1101" => d <= "00110110"; -- ..##.##.
                when x"cc" & "1110" => d <= "00110110"; -- ..##.##.
                when x"cc" & "1111" => d <= "00110110"; -- ..##.##.

                when x"cd" & "0000" => d <= "00000000"; -- ........
                when x"cd" & "0001" => d <= "00000000"; -- ........
                when x"cd" & "0010" => d <= "00000000"; -- ........
                when x"cd" & "0011" => d <= "00000000"; -- ........
                when x"cd" & "0100" => d <= "00000000"; -- ........
                when x"cd" & "0101" => d <= "11111111"; -- ########
                when x"cd" & "0110" => d <= "00000000"; -- ........
                when x"cd" & "0111" => d <= "11111111"; -- ########
                when x"cd" & "1000" => d <= "00000000"; -- ........
                when x"cd" & "1001" => d <= "00000000"; -- ........
                when x"cd" & "1010" => d <= "00000000"; -- ........
                when x"cd" & "1011" => d <= "00000000"; -- ........
                when x"cd" & "1100" => d <= "00000000"; -- ........
                when x"cd" & "1101" => d <= "00000000"; -- ........
                when x"cd" & "1110" => d <= "00000000"; -- ........
                when x"cd" & "1111" => d <= "00000000"; -- ........

                when x"ce" & "0000" => d <= "00110110"; -- ..##.##.
                when x"ce" & "0001" => d <= "00110110"; -- ..##.##.
                when x"ce" & "0010" => d <= "00110110"; -- ..##.##.
                when x"ce" & "0011" => d <= "00110110"; -- ..##.##.
                when x"ce" & "0100" => d <= "00110110"; -- ..##.##.
                when x"ce" & "0101" => d <= "11110111"; -- ####.###
                when x"ce" & "0110" => d <= "00000000"; -- ........
                when x"ce" & "0111" => d <= "11110111"; -- ####.###
                when x"ce" & "1000" => d <= "00110110"; -- ..##.##.
                when x"ce" & "1001" => d <= "00110110"; -- ..##.##.
                when x"ce" & "1010" => d <= "00110110"; -- ..##.##.
                when x"ce" & "1011" => d <= "00110110"; -- ..##.##.
                when x"ce" & "1100" => d <= "00110110"; -- ..##.##.
                when x"ce" & "1101" => d <= "00110110"; -- ..##.##.
                when x"ce" & "1110" => d <= "00110110"; -- ..##.##.
                when x"ce" & "1111" => d <= "00110110"; -- ..##.##.

                when x"cf" & "0000" => d <= "00011000"; -- ...##...
                when x"cf" & "0001" => d <= "00011000"; -- ...##...
                when x"cf" & "0010" => d <= "00011000"; -- ...##...
                when x"cf" & "0011" => d <= "00011000"; -- ...##...
                when x"cf" & "0100" => d <= "00011000"; -- ...##...
                when x"cf" & "0101" => d <= "11111111"; -- ########
                when x"cf" & "0110" => d <= "00000000"; -- ........
                when x"cf" & "0111" => d <= "11111111"; -- ########
                when x"cf" & "1000" => d <= "00000000"; -- ........
                when x"cf" & "1001" => d <= "00000000"; -- ........
                when x"cf" & "1010" => d <= "00000000"; -- ........
                when x"cf" & "1011" => d <= "00000000"; -- ........
                when x"cf" & "1100" => d <= "00000000"; -- ........
                when x"cf" & "1101" => d <= "00000000"; -- ........
                when x"cf" & "1110" => d <= "00000000"; -- ........
                when x"cf" & "1111" => d <= "00000000"; -- ........

                when x"d0" & "0000" => d <= "00110110"; -- ..##.##.
                when x"d0" & "0001" => d <= "00110110"; -- ..##.##.
                when x"d0" & "0010" => d <= "00110110"; -- ..##.##.
                when x"d0" & "0011" => d <= "00110110"; -- ..##.##.
                when x"d0" & "0100" => d <= "00110110"; -- ..##.##.
                when x"d0" & "0101" => d <= "00110110"; -- ..##.##.
                when x"d0" & "0110" => d <= "00110110"; -- ..##.##.
                when x"d0" & "0111" => d <= "11111111"; -- ########
                when x"d0" & "1000" => d <= "00000000"; -- ........
                when x"d0" & "1001" => d <= "00000000"; -- ........
                when x"d0" & "1010" => d <= "00000000"; -- ........
                when x"d0" & "1011" => d <= "00000000"; -- ........
                when x"d0" & "1100" => d <= "00000000"; -- ........
                when x"d0" & "1101" => d <= "00000000"; -- ........
                when x"d0" & "1110" => d <= "00000000"; -- ........
                when x"d0" & "1111" => d <= "00000000"; -- ........

                when x"d1" & "0000" => d <= "00000000"; -- ........
                when x"d1" & "0001" => d <= "00000000"; -- ........
                when x"d1" & "0010" => d <= "00000000"; -- ........
                when x"d1" & "0011" => d <= "00000000"; -- ........
                when x"d1" & "0100" => d <= "00000000"; -- ........
                when x"d1" & "0101" => d <= "11111111"; -- ########
                when x"d1" & "0110" => d <= "00000000"; -- ........
                when x"d1" & "0111" => d <= "11111111"; -- ########
                when x"d1" & "1000" => d <= "00011000"; -- ...##...
                when x"d1" & "1001" => d <= "00011000"; -- ...##...
                when x"d1" & "1010" => d <= "00011000"; -- ...##...
                when x"d1" & "1011" => d <= "00011000"; -- ...##...
                when x"d1" & "1100" => d <= "00011000"; -- ...##...
                when x"d1" & "1101" => d <= "00011000"; -- ...##...
                when x"d1" & "1110" => d <= "00011000"; -- ...##...
                when x"d1" & "1111" => d <= "00011000"; -- ...##...

                when x"d2" & "0000" => d <= "00000000"; -- ........
                when x"d2" & "0001" => d <= "00000000"; -- ........
                when x"d2" & "0010" => d <= "00000000"; -- ........
                when x"d2" & "0011" => d <= "00000000"; -- ........
                when x"d2" & "0100" => d <= "00000000"; -- ........
                when x"d2" & "0101" => d <= "00000000"; -- ........
                when x"d2" & "0110" => d <= "00000000"; -- ........
                when x"d2" & "0111" => d <= "11111111"; -- ########
                when x"d2" & "1000" => d <= "00110110"; -- ..##.##.
                when x"d2" & "1001" => d <= "00110110"; -- ..##.##.
                when x"d2" & "1010" => d <= "00110110"; -- ..##.##.
                when x"d2" & "1011" => d <= "00110110"; -- ..##.##.
                when x"d2" & "1100" => d <= "00110110"; -- ..##.##.
                when x"d2" & "1101" => d <= "00110110"; -- ..##.##.
                when x"d2" & "1110" => d <= "00110110"; -- ..##.##.
                when x"d2" & "1111" => d <= "00110110"; -- ..##.##.

                when x"d3" & "0000" => d <= "00110110"; -- ..##.##.
                when x"d3" & "0001" => d <= "00110110"; -- ..##.##.
                when x"d3" & "0010" => d <= "00110110"; -- ..##.##.
                when x"d3" & "0011" => d <= "00110110"; -- ..##.##.
                when x"d3" & "0100" => d <= "00110110"; -- ..##.##.
                when x"d3" & "0101" => d <= "00110110"; -- ..##.##.
                when x"d3" & "0110" => d <= "00110110"; -- ..##.##.
                when x"d3" & "0111" => d <= "00111111"; -- ..######
                when x"d3" & "1000" => d <= "00000000"; -- ........
                when x"d3" & "1001" => d <= "00000000"; -- ........
                when x"d3" & "1010" => d <= "00000000"; -- ........
                when x"d3" & "1011" => d <= "00000000"; -- ........
                when x"d3" & "1100" => d <= "00000000"; -- ........
                when x"d3" & "1101" => d <= "00000000"; -- ........
                when x"d3" & "1110" => d <= "00000000"; -- ........
                when x"d3" & "1111" => d <= "00000000"; -- ........

                when x"d4" & "0000" => d <= "00011000"; -- ...##...
                when x"d4" & "0001" => d <= "00011000"; -- ...##...
                when x"d4" & "0010" => d <= "00011000"; -- ...##...
                when x"d4" & "0011" => d <= "00011000"; -- ...##...
                when x"d4" & "0100" => d <= "00011000"; -- ...##...
                when x"d4" & "0101" => d <= "00011111"; -- ...#####
                when x"d4" & "0110" => d <= "00011000"; -- ...##...
                when x"d4" & "0111" => d <= "00011111"; -- ...#####
                when x"d4" & "1000" => d <= "00000000"; -- ........
                when x"d4" & "1001" => d <= "00000000"; -- ........
                when x"d4" & "1010" => d <= "00000000"; -- ........
                when x"d4" & "1011" => d <= "00000000"; -- ........
                when x"d4" & "1100" => d <= "00000000"; -- ........
                when x"d4" & "1101" => d <= "00000000"; -- ........
                when x"d4" & "1110" => d <= "00000000"; -- ........
                when x"d4" & "1111" => d <= "00000000"; -- ........

                when x"d5" & "0000" => d <= "00000000"; -- ........
                when x"d5" & "0001" => d <= "00000000"; -- ........
                when x"d5" & "0010" => d <= "00000000"; -- ........
                when x"d5" & "0011" => d <= "00000000"; -- ........
                when x"d5" & "0100" => d <= "00000000"; -- ........
                when x"d5" & "0101" => d <= "00011111"; -- ...#####
                when x"d5" & "0110" => d <= "00011000"; -- ...##...
                when x"d5" & "0111" => d <= "00011111"; -- ...#####
                when x"d5" & "1000" => d <= "00011000"; -- ...##...
                when x"d5" & "1001" => d <= "00011000"; -- ...##...
                when x"d5" & "1010" => d <= "00011000"; -- ...##...
                when x"d5" & "1011" => d <= "00011000"; -- ...##...
                when x"d5" & "1100" => d <= "00011000"; -- ...##...
                when x"d5" & "1101" => d <= "00011000"; -- ...##...
                when x"d5" & "1110" => d <= "00011000"; -- ...##...
                when x"d5" & "1111" => d <= "00011000"; -- ...##...

                when x"d6" & "0000" => d <= "00000000"; -- ........
                when x"d6" & "0001" => d <= "00000000"; -- ........
                when x"d6" & "0010" => d <= "00000000"; -- ........
                when x"d6" & "0011" => d <= "00000000"; -- ........
                when x"d6" & "0100" => d <= "00000000"; -- ........
                when x"d6" & "0101" => d <= "00000000"; -- ........
                when x"d6" & "0110" => d <= "00000000"; -- ........
                when x"d6" & "0111" => d <= "00111111"; -- ..######
                when x"d6" & "1000" => d <= "00110110"; -- ..##.##.
                when x"d6" & "1001" => d <= "00110110"; -- ..##.##.
                when x"d6" & "1010" => d <= "00110110"; -- ..##.##.
                when x"d6" & "1011" => d <= "00110110"; -- ..##.##.
                when x"d6" & "1100" => d <= "00110110"; -- ..##.##.
                when x"d6" & "1101" => d <= "00110110"; -- ..##.##.
                when x"d6" & "1110" => d <= "00110110"; -- ..##.##.
                when x"d6" & "1111" => d <= "00110110"; -- ..##.##.

                when x"d7" & "0000" => d <= "00110110"; -- ..##.##.
                when x"d7" & "0001" => d <= "00110110"; -- ..##.##.
                when x"d7" & "0010" => d <= "00110110"; -- ..##.##.
                when x"d7" & "0011" => d <= "00110110"; -- ..##.##.
                when x"d7" & "0100" => d <= "00110110"; -- ..##.##.
                when x"d7" & "0101" => d <= "00110110"; -- ..##.##.
                when x"d7" & "0110" => d <= "00110110"; -- ..##.##.
                when x"d7" & "0111" => d <= "11111111"; -- ########
                when x"d7" & "1000" => d <= "00110110"; -- ..##.##.
                when x"d7" & "1001" => d <= "00110110"; -- ..##.##.
                when x"d7" & "1010" => d <= "00110110"; -- ..##.##.
                when x"d7" & "1011" => d <= "00110110"; -- ..##.##.
                when x"d7" & "1100" => d <= "00110110"; -- ..##.##.
                when x"d7" & "1101" => d <= "00110110"; -- ..##.##.
                when x"d7" & "1110" => d <= "00110110"; -- ..##.##.
                when x"d7" & "1111" => d <= "00110110"; -- ..##.##.

                when x"d8" & "0000" => d <= "00011000"; -- ...##...
                when x"d8" & "0001" => d <= "00011000"; -- ...##...
                when x"d8" & "0010" => d <= "00011000"; -- ...##...
                when x"d8" & "0011" => d <= "00011000"; -- ...##...
                when x"d8" & "0100" => d <= "00011000"; -- ...##...
                when x"d8" & "0101" => d <= "11111111"; -- ########
                when x"d8" & "0110" => d <= "00011000"; -- ...##...
                when x"d8" & "0111" => d <= "11111111"; -- ########
                when x"d8" & "1000" => d <= "00011000"; -- ...##...
                when x"d8" & "1001" => d <= "00011000"; -- ...##...
                when x"d8" & "1010" => d <= "00011000"; -- ...##...
                when x"d8" & "1011" => d <= "00011000"; -- ...##...
                when x"d8" & "1100" => d <= "00011000"; -- ...##...
                when x"d8" & "1101" => d <= "00011000"; -- ...##...
                when x"d8" & "1110" => d <= "00011000"; -- ...##...
                when x"d8" & "1111" => d <= "00011000"; -- ...##...

                when x"d9" & "0000" => d <= "00011000"; -- ...##...
                when x"d9" & "0001" => d <= "00011000"; -- ...##...
                when x"d9" & "0010" => d <= "00011000"; -- ...##...
                when x"d9" & "0011" => d <= "00011000"; -- ...##...
                when x"d9" & "0100" => d <= "00011000"; -- ...##...
                when x"d9" & "0101" => d <= "00011000"; -- ...##...
                when x"d9" & "0110" => d <= "00011000"; -- ...##...
                when x"d9" & "0111" => d <= "11111000"; -- #####...
                when x"d9" & "1000" => d <= "00000000"; -- ........
                when x"d9" & "1001" => d <= "00000000"; -- ........
                when x"d9" & "1010" => d <= "00000000"; -- ........
                when x"d9" & "1011" => d <= "00000000"; -- ........
                when x"d9" & "1100" => d <= "00000000"; -- ........
                when x"d9" & "1101" => d <= "00000000"; -- ........
                when x"d9" & "1110" => d <= "00000000"; -- ........
                when x"d9" & "1111" => d <= "00000000"; -- ........

                when x"da" & "0000" => d <= "00000000"; -- ........
                when x"da" & "0001" => d <= "00000000"; -- ........
                when x"da" & "0010" => d <= "00000000"; -- ........
                when x"da" & "0011" => d <= "00000000"; -- ........
                when x"da" & "0100" => d <= "00000000"; -- ........
                when x"da" & "0101" => d <= "00000000"; -- ........
                when x"da" & "0110" => d <= "00000000"; -- ........
                when x"da" & "0111" => d <= "00011111"; -- ...#####
                when x"da" & "1000" => d <= "00011000"; -- ...##...
                when x"da" & "1001" => d <= "00011000"; -- ...##...
                when x"da" & "1010" => d <= "00011000"; -- ...##...
                when x"da" & "1011" => d <= "00011000"; -- ...##...
                when x"da" & "1100" => d <= "00011000"; -- ...##...
                when x"da" & "1101" => d <= "00011000"; -- ...##...
                when x"da" & "1110" => d <= "00011000"; -- ...##...
                when x"da" & "1111" => d <= "00011000"; -- ...##...

                when x"db" & "0000" => d <= "11111111"; -- ########
                when x"db" & "0001" => d <= "11111111"; -- ########
                when x"db" & "0010" => d <= "11111111"; -- ########
                when x"db" & "0011" => d <= "11111111"; -- ########
                when x"db" & "0100" => d <= "11111111"; -- ########
                when x"db" & "0101" => d <= "11111111"; -- ########
                when x"db" & "0110" => d <= "11111111"; -- ########
                when x"db" & "0111" => d <= "11111111"; -- ########
                when x"db" & "1000" => d <= "11111111"; -- ########
                when x"db" & "1001" => d <= "11111111"; -- ########
                when x"db" & "1010" => d <= "11111111"; -- ########
                when x"db" & "1011" => d <= "11111111"; -- ########
                when x"db" & "1100" => d <= "11111111"; -- ########
                when x"db" & "1101" => d <= "11111111"; -- ########
                when x"db" & "1110" => d <= "11111111"; -- ########
                when x"db" & "1111" => d <= "11111111"; -- ########

                when x"dc" & "0000" => d <= "00000000"; -- ........
                when x"dc" & "0001" => d <= "00000000"; -- ........
                when x"dc" & "0010" => d <= "00000000"; -- ........
                when x"dc" & "0011" => d <= "00000000"; -- ........
                when x"dc" & "0100" => d <= "00000000"; -- ........
                when x"dc" & "0101" => d <= "00000000"; -- ........
                when x"dc" & "0110" => d <= "00000000"; -- ........
                when x"dc" & "0111" => d <= "11111111"; -- ########
                when x"dc" & "1000" => d <= "11111111"; -- ########
                when x"dc" & "1001" => d <= "11111111"; -- ########
                when x"dc" & "1010" => d <= "11111111"; -- ########
                when x"dc" & "1011" => d <= "11111111"; -- ########
                when x"dc" & "1100" => d <= "11111111"; -- ########
                when x"dc" & "1101" => d <= "11111111"; -- ########
                when x"dc" & "1110" => d <= "11111111"; -- ########
                when x"dc" & "1111" => d <= "11111111"; -- ########

                when x"dd" & "0000" => d <= "11110000"; -- ####....
                when x"dd" & "0001" => d <= "11110000"; -- ####....
                when x"dd" & "0010" => d <= "11110000"; -- ####....
                when x"dd" & "0011" => d <= "11110000"; -- ####....
                when x"dd" & "0100" => d <= "11110000"; -- ####....
                when x"dd" & "0101" => d <= "11110000"; -- ####....
                when x"dd" & "0110" => d <= "11110000"; -- ####....
                when x"dd" & "0111" => d <= "11110000"; -- ####....
                when x"dd" & "1000" => d <= "11110000"; -- ####....
                when x"dd" & "1001" => d <= "11110000"; -- ####....
                when x"dd" & "1010" => d <= "11110000"; -- ####....
                when x"dd" & "1011" => d <= "11110000"; -- ####....
                when x"dd" & "1100" => d <= "11110000"; -- ####....
                when x"dd" & "1101" => d <= "11110000"; -- ####....
                when x"dd" & "1110" => d <= "11110000"; -- ####....
                when x"dd" & "1111" => d <= "11110000"; -- ####....

                when x"de" & "0000" => d <= "00001111"; -- ....####
                when x"de" & "0001" => d <= "00001111"; -- ....####
                when x"de" & "0010" => d <= "00001111"; -- ....####
                when x"de" & "0011" => d <= "00001111"; -- ....####
                when x"de" & "0100" => d <= "00001111"; -- ....####
                when x"de" & "0101" => d <= "00001111"; -- ....####
                when x"de" & "0110" => d <= "00001111"; -- ....####
                when x"de" & "0111" => d <= "00001111"; -- ....####
                when x"de" & "1000" => d <= "00001111"; -- ....####
                when x"de" & "1001" => d <= "00001111"; -- ....####
                when x"de" & "1010" => d <= "00001111"; -- ....####
                when x"de" & "1011" => d <= "00001111"; -- ....####
                when x"de" & "1100" => d <= "00001111"; -- ....####
                when x"de" & "1101" => d <= "00001111"; -- ....####
                when x"de" & "1110" => d <= "00001111"; -- ....####
                when x"de" & "1111" => d <= "00001111"; -- ....####

                when x"df" & "0000" => d <= "11111111"; -- ########
                when x"df" & "0001" => d <= "11111111"; -- ########
                when x"df" & "0010" => d <= "11111111"; -- ########
                when x"df" & "0011" => d <= "11111111"; -- ########
                when x"df" & "0100" => d <= "11111111"; -- ########
                when x"df" & "0101" => d <= "11111111"; -- ########
                when x"df" & "0110" => d <= "11111111"; -- ########
                when x"df" & "0111" => d <= "00000000"; -- ........
                when x"df" & "1000" => d <= "00000000"; -- ........
                when x"df" & "1001" => d <= "00000000"; -- ........
                when x"df" & "1010" => d <= "00000000"; -- ........
                when x"df" & "1011" => d <= "00000000"; -- ........
                when x"df" & "1100" => d <= "00000000"; -- ........
                when x"df" & "1101" => d <= "00000000"; -- ........
                when x"df" & "1110" => d <= "00000000"; -- ........
                when x"df" & "1111" => d <= "00000000"; -- ........

                when x"e0" & "0000" => d <= "00000000"; -- ........
                when x"e0" & "0001" => d <= "00000000"; -- ........
                when x"e0" & "0010" => d <= "00000000"; -- ........
                when x"e0" & "0011" => d <= "00000000"; -- ........
                when x"e0" & "0100" => d <= "00000000"; -- ........
                when x"e0" & "0101" => d <= "01110110"; -- .###.##.
                when x"e0" & "0110" => d <= "11011100"; -- ##.###..
                when x"e0" & "0111" => d <= "11011000"; -- ##.##...
                when x"e0" & "1000" => d <= "11011000"; -- ##.##...
                when x"e0" & "1001" => d <= "11011000"; -- ##.##...
                when x"e0" & "1010" => d <= "11011100"; -- ##.###..
                when x"e0" & "1011" => d <= "01110110"; -- .###.##.
                when x"e0" & "1100" => d <= "00000000"; -- ........
                when x"e0" & "1101" => d <= "00000000"; -- ........
                when x"e0" & "1110" => d <= "00000000"; -- ........
                when x"e0" & "1111" => d <= "00000000"; -- ........

                when x"e1" & "0000" => d <= "00000000"; -- ........
                when x"e1" & "0001" => d <= "00000000"; -- ........
                when x"e1" & "0010" => d <= "01111000"; -- .####...
                when x"e1" & "0011" => d <= "11001100"; -- ##..##..
                when x"e1" & "0100" => d <= "11001100"; -- ##..##..
                when x"e1" & "0101" => d <= "11001100"; -- ##..##..
                when x"e1" & "0110" => d <= "11011000"; -- ##.##...
                when x"e1" & "0111" => d <= "11001100"; -- ##..##..
                when x"e1" & "1000" => d <= "11000110"; -- ##...##.
                when x"e1" & "1001" => d <= "11000110"; -- ##...##.
                when x"e1" & "1010" => d <= "11000110"; -- ##...##.
                when x"e1" & "1011" => d <= "11001100"; -- ##..##..
                when x"e1" & "1100" => d <= "00000000"; -- ........
                when x"e1" & "1101" => d <= "00000000"; -- ........
                when x"e1" & "1110" => d <= "00000000"; -- ........
                when x"e1" & "1111" => d <= "00000000"; -- ........

                when x"e2" & "0000" => d <= "00000000"; -- ........
                when x"e2" & "0001" => d <= "00000000"; -- ........
                when x"e2" & "0010" => d <= "11111110"; -- #######.
                when x"e2" & "0011" => d <= "11000110"; -- ##...##.
                when x"e2" & "0100" => d <= "11000110"; -- ##...##.
                when x"e2" & "0101" => d <= "11000000"; -- ##......
                when x"e2" & "0110" => d <= "11000000"; -- ##......
                when x"e2" & "0111" => d <= "11000000"; -- ##......
                when x"e2" & "1000" => d <= "11000000"; -- ##......
                when x"e2" & "1001" => d <= "11000000"; -- ##......
                when x"e2" & "1010" => d <= "11000000"; -- ##......
                when x"e2" & "1011" => d <= "11000000"; -- ##......
                when x"e2" & "1100" => d <= "00000000"; -- ........
                when x"e2" & "1101" => d <= "00000000"; -- ........
                when x"e2" & "1110" => d <= "00000000"; -- ........
                when x"e2" & "1111" => d <= "00000000"; -- ........

                when x"e3" & "0000" => d <= "00000000"; -- ........
                when x"e3" & "0001" => d <= "00000000"; -- ........
                when x"e3" & "0010" => d <= "00000000"; -- ........
                when x"e3" & "0011" => d <= "00000000"; -- ........
                when x"e3" & "0100" => d <= "11111110"; -- #######.
                when x"e3" & "0101" => d <= "01101100"; -- .##.##..
                when x"e3" & "0110" => d <= "01101100"; -- .##.##..
                when x"e3" & "0111" => d <= "01101100"; -- .##.##..
                when x"e3" & "1000" => d <= "01101100"; -- .##.##..
                when x"e3" & "1001" => d <= "01101100"; -- .##.##..
                when x"e3" & "1010" => d <= "01101100"; -- .##.##..
                when x"e3" & "1011" => d <= "01101100"; -- .##.##..
                when x"e3" & "1100" => d <= "00000000"; -- ........
                when x"e3" & "1101" => d <= "00000000"; -- ........
                when x"e3" & "1110" => d <= "00000000"; -- ........
                when x"e3" & "1111" => d <= "00000000"; -- ........

                when x"e4" & "0000" => d <= "00000000"; -- ........
                when x"e4" & "0001" => d <= "00000000"; -- ........
                when x"e4" & "0010" => d <= "00000000"; -- ........
                when x"e4" & "0011" => d <= "11111110"; -- #######.
                when x"e4" & "0100" => d <= "11000110"; -- ##...##.
                when x"e4" & "0101" => d <= "01100000"; -- .##.....
                when x"e4" & "0110" => d <= "00110000"; -- ..##....
                when x"e4" & "0111" => d <= "00011000"; -- ...##...
                when x"e4" & "1000" => d <= "00110000"; -- ..##....
                when x"e4" & "1001" => d <= "01100000"; -- .##.....
                when x"e4" & "1010" => d <= "11000110"; -- ##...##.
                when x"e4" & "1011" => d <= "11111110"; -- #######.
                when x"e4" & "1100" => d <= "00000000"; -- ........
                when x"e4" & "1101" => d <= "00000000"; -- ........
                when x"e4" & "1110" => d <= "00000000"; -- ........
                when x"e4" & "1111" => d <= "00000000"; -- ........

                when x"e5" & "0000" => d <= "00000000"; -- ........
                when x"e5" & "0001" => d <= "00000000"; -- ........
                when x"e5" & "0010" => d <= "00000000"; -- ........
                when x"e5" & "0011" => d <= "00000000"; -- ........
                when x"e5" & "0100" => d <= "00000000"; -- ........
                when x"e5" & "0101" => d <= "01111110"; -- .######.
                when x"e5" & "0110" => d <= "11011000"; -- ##.##...
                when x"e5" & "0111" => d <= "11011000"; -- ##.##...
                when x"e5" & "1000" => d <= "11011000"; -- ##.##...
                when x"e5" & "1001" => d <= "11011000"; -- ##.##...
                when x"e5" & "1010" => d <= "11011000"; -- ##.##...
                when x"e5" & "1011" => d <= "01110000"; -- .###....
                when x"e5" & "1100" => d <= "00000000"; -- ........
                when x"e5" & "1101" => d <= "00000000"; -- ........
                when x"e5" & "1110" => d <= "00000000"; -- ........
                when x"e5" & "1111" => d <= "00000000"; -- ........

                when x"e6" & "0000" => d <= "00000000"; -- ........
                when x"e6" & "0001" => d <= "00000000"; -- ........
                when x"e6" & "0010" => d <= "00000000"; -- ........
                when x"e6" & "0011" => d <= "00000000"; -- ........
                when x"e6" & "0100" => d <= "01100110"; -- .##..##.
                when x"e6" & "0101" => d <= "01100110"; -- .##..##.
                when x"e6" & "0110" => d <= "01100110"; -- .##..##.
                when x"e6" & "0111" => d <= "01100110"; -- .##..##.
                when x"e6" & "1000" => d <= "01100110"; -- .##..##.
                when x"e6" & "1001" => d <= "01111100"; -- .#####..
                when x"e6" & "1010" => d <= "01100000"; -- .##.....
                when x"e6" & "1011" => d <= "01100000"; -- .##.....
                when x"e6" & "1100" => d <= "11000000"; -- ##......
                when x"e6" & "1101" => d <= "00000000"; -- ........
                when x"e6" & "1110" => d <= "00000000"; -- ........
                when x"e6" & "1111" => d <= "00000000"; -- ........

                when x"e7" & "0000" => d <= "00000000"; -- ........
                when x"e7" & "0001" => d <= "00000000"; -- ........
                when x"e7" & "0010" => d <= "00000000"; -- ........
                when x"e7" & "0011" => d <= "00000000"; -- ........
                when x"e7" & "0100" => d <= "01110110"; -- .###.##.
                when x"e7" & "0101" => d <= "11011100"; -- ##.###..
                when x"e7" & "0110" => d <= "00011000"; -- ...##...
                when x"e7" & "0111" => d <= "00011000"; -- ...##...
                when x"e7" & "1000" => d <= "00011000"; -- ...##...
                when x"e7" & "1001" => d <= "00011000"; -- ...##...
                when x"e7" & "1010" => d <= "00011000"; -- ...##...
                when x"e7" & "1011" => d <= "00011000"; -- ...##...
                when x"e7" & "1100" => d <= "00000000"; -- ........
                when x"e7" & "1101" => d <= "00000000"; -- ........
                when x"e7" & "1110" => d <= "00000000"; -- ........
                when x"e7" & "1111" => d <= "00000000"; -- ........

                when x"e8" & "0000" => d <= "00000000"; -- ........
                when x"e8" & "0001" => d <= "00000000"; -- ........
                when x"e8" & "0010" => d <= "00000000"; -- ........
                when x"e8" & "0011" => d <= "01111110"; -- .######.
                when x"e8" & "0100" => d <= "00011000"; -- ...##...
                when x"e8" & "0101" => d <= "00111100"; -- ..####..
                when x"e8" & "0110" => d <= "01100110"; -- .##..##.
                when x"e8" & "0111" => d <= "01100110"; -- .##..##.
                when x"e8" & "1000" => d <= "01100110"; -- .##..##.
                when x"e8" & "1001" => d <= "00111100"; -- ..####..
                when x"e8" & "1010" => d <= "00011000"; -- ...##...
                when x"e8" & "1011" => d <= "01111110"; -- .######.
                when x"e8" & "1100" => d <= "00000000"; -- ........
                when x"e8" & "1101" => d <= "00000000"; -- ........
                when x"e8" & "1110" => d <= "00000000"; -- ........
                when x"e8" & "1111" => d <= "00000000"; -- ........

                when x"e9" & "0000" => d <= "00000000"; -- ........
                when x"e9" & "0001" => d <= "00000000"; -- ........
                when x"e9" & "0010" => d <= "00000000"; -- ........
                when x"e9" & "0011" => d <= "00111000"; -- ..###...
                when x"e9" & "0100" => d <= "01101100"; -- .##.##..
                when x"e9" & "0101" => d <= "11000110"; -- ##...##.
                when x"e9" & "0110" => d <= "11000110"; -- ##...##.
                when x"e9" & "0111" => d <= "11111110"; -- #######.
                when x"e9" & "1000" => d <= "11000110"; -- ##...##.
                when x"e9" & "1001" => d <= "11000110"; -- ##...##.
                when x"e9" & "1010" => d <= "01101100"; -- .##.##..
                when x"e9" & "1011" => d <= "00111000"; -- ..###...
                when x"e9" & "1100" => d <= "00000000"; -- ........
                when x"e9" & "1101" => d <= "00000000"; -- ........
                when x"e9" & "1110" => d <= "00000000"; -- ........
                when x"e9" & "1111" => d <= "00000000"; -- ........

                when x"ea" & "0000" => d <= "00000000"; -- ........
                when x"ea" & "0001" => d <= "00000000"; -- ........
                when x"ea" & "0010" => d <= "00111000"; -- ..###...
                when x"ea" & "0011" => d <= "01101100"; -- .##.##..
                when x"ea" & "0100" => d <= "11000110"; -- ##...##.
                when x"ea" & "0101" => d <= "11000110"; -- ##...##.
                when x"ea" & "0110" => d <= "11000110"; -- ##...##.
                when x"ea" & "0111" => d <= "01101100"; -- .##.##..
                when x"ea" & "1000" => d <= "01101100"; -- .##.##..
                when x"ea" & "1001" => d <= "01101100"; -- .##.##..
                when x"ea" & "1010" => d <= "01101100"; -- .##.##..
                when x"ea" & "1011" => d <= "11101110"; -- ###.###.
                when x"ea" & "1100" => d <= "00000000"; -- ........
                when x"ea" & "1101" => d <= "00000000"; -- ........
                when x"ea" & "1110" => d <= "00000000"; -- ........
                when x"ea" & "1111" => d <= "00000000"; -- ........

                when x"eb" & "0000" => d <= "00000000"; -- ........
                when x"eb" & "0001" => d <= "00000000"; -- ........
                when x"eb" & "0010" => d <= "00011110"; -- ...####.
                when x"eb" & "0011" => d <= "00110000"; -- ..##....
                when x"eb" & "0100" => d <= "00011000"; -- ...##...
                when x"eb" & "0101" => d <= "00001100"; -- ....##..
                when x"eb" & "0110" => d <= "00111110"; -- ..#####.
                when x"eb" & "0111" => d <= "01100110"; -- .##..##.
                when x"eb" & "1000" => d <= "01100110"; -- .##..##.
                when x"eb" & "1001" => d <= "01100110"; -- .##..##.
                when x"eb" & "1010" => d <= "01100110"; -- .##..##.
                when x"eb" & "1011" => d <= "00111100"; -- ..####..
                when x"eb" & "1100" => d <= "00000000"; -- ........
                when x"eb" & "1101" => d <= "00000000"; -- ........
                when x"eb" & "1110" => d <= "00000000"; -- ........
                when x"eb" & "1111" => d <= "00000000"; -- ........

                when x"ec" & "0000" => d <= "00000000"; -- ........
                when x"ec" & "0001" => d <= "00000000"; -- ........
                when x"ec" & "0010" => d <= "00000000"; -- ........
                when x"ec" & "0011" => d <= "00000000"; -- ........
                when x"ec" & "0100" => d <= "00000000"; -- ........
                when x"ec" & "0101" => d <= "01111110"; -- .######.
                when x"ec" & "0110" => d <= "11011011"; -- ##.##.##
                when x"ec" & "0111" => d <= "11011011"; -- ##.##.##
                when x"ec" & "1000" => d <= "11011011"; -- ##.##.##
                when x"ec" & "1001" => d <= "01111110"; -- .######.
                when x"ec" & "1010" => d <= "00000000"; -- ........
                when x"ec" & "1011" => d <= "00000000"; -- ........
                when x"ec" & "1100" => d <= "00000000"; -- ........
                when x"ec" & "1101" => d <= "00000000"; -- ........
                when x"ec" & "1110" => d <= "00000000"; -- ........
                when x"ec" & "1111" => d <= "00000000"; -- ........

                when x"ed" & "0000" => d <= "00000000"; -- ........
                when x"ed" & "0001" => d <= "00000000"; -- ........
                when x"ed" & "0010" => d <= "00000000"; -- ........
                when x"ed" & "0011" => d <= "00000011"; -- ......##
                when x"ed" & "0100" => d <= "00000110"; -- .....##.
                when x"ed" & "0101" => d <= "01111110"; -- .######.
                when x"ed" & "0110" => d <= "11011011"; -- ##.##.##
                when x"ed" & "0111" => d <= "11011011"; -- ##.##.##
                when x"ed" & "1000" => d <= "11110011"; -- ####..##
                when x"ed" & "1001" => d <= "01111110"; -- .######.
                when x"ed" & "1010" => d <= "01100000"; -- .##.....
                when x"ed" & "1011" => d <= "11000000"; -- ##......
                when x"ed" & "1100" => d <= "00000000"; -- ........
                when x"ed" & "1101" => d <= "00000000"; -- ........
                when x"ed" & "1110" => d <= "00000000"; -- ........
                when x"ed" & "1111" => d <= "00000000"; -- ........

                when x"ee" & "0000" => d <= "00000000"; -- ........
                when x"ee" & "0001" => d <= "00000000"; -- ........
                when x"ee" & "0010" => d <= "00011100"; -- ...###..
                when x"ee" & "0011" => d <= "00110000"; -- ..##....
                when x"ee" & "0100" => d <= "01100000"; -- .##.....
                when x"ee" & "0101" => d <= "01100000"; -- .##.....
                when x"ee" & "0110" => d <= "01111100"; -- .#####..
                when x"ee" & "0111" => d <= "01100000"; -- .##.....
                when x"ee" & "1000" => d <= "01100000"; -- .##.....
                when x"ee" & "1001" => d <= "01100000"; -- .##.....
                when x"ee" & "1010" => d <= "00110000"; -- ..##....
                when x"ee" & "1011" => d <= "00011100"; -- ...###..
                when x"ee" & "1100" => d <= "00000000"; -- ........
                when x"ee" & "1101" => d <= "00000000"; -- ........
                when x"ee" & "1110" => d <= "00000000"; -- ........
                when x"ee" & "1111" => d <= "00000000"; -- ........

                when x"ef" & "0000" => d <= "00000000"; -- ........
                when x"ef" & "0001" => d <= "00000000"; -- ........
                when x"ef" & "0010" => d <= "00000000"; -- ........
                when x"ef" & "0011" => d <= "01111100"; -- .#####..
                when x"ef" & "0100" => d <= "11000110"; -- ##...##.
                when x"ef" & "0101" => d <= "11000110"; -- ##...##.
                when x"ef" & "0110" => d <= "11000110"; -- ##...##.
                when x"ef" & "0111" => d <= "11000110"; -- ##...##.
                when x"ef" & "1000" => d <= "11000110"; -- ##...##.
                when x"ef" & "1001" => d <= "11000110"; -- ##...##.
                when x"ef" & "1010" => d <= "11000110"; -- ##...##.
                when x"ef" & "1011" => d <= "11000110"; -- ##...##.
                when x"ef" & "1100" => d <= "00000000"; -- ........
                when x"ef" & "1101" => d <= "00000000"; -- ........
                when x"ef" & "1110" => d <= "00000000"; -- ........
                when x"ef" & "1111" => d <= "00000000"; -- ........

                when x"f0" & "0000" => d <= "00000000"; -- ........
                when x"f0" & "0001" => d <= "00000000"; -- ........
                when x"f0" & "0010" => d <= "00000000"; -- ........
                when x"f0" & "0011" => d <= "00000000"; -- ........
                when x"f0" & "0100" => d <= "11111110"; -- #######.
                when x"f0" & "0101" => d <= "00000000"; -- ........
                when x"f0" & "0110" => d <= "00000000"; -- ........
                when x"f0" & "0111" => d <= "11111110"; -- #######.
                when x"f0" & "1000" => d <= "00000000"; -- ........
                when x"f0" & "1001" => d <= "00000000"; -- ........
                when x"f0" & "1010" => d <= "11111110"; -- #######.
                when x"f0" & "1011" => d <= "00000000"; -- ........
                when x"f0" & "1100" => d <= "00000000"; -- ........
                when x"f0" & "1101" => d <= "00000000"; -- ........
                when x"f0" & "1110" => d <= "00000000"; -- ........
                when x"f0" & "1111" => d <= "00000000"; -- ........

                when x"f1" & "0000" => d <= "00000000"; -- ........
                when x"f1" & "0001" => d <= "00000000"; -- ........
                when x"f1" & "0010" => d <= "00000000"; -- ........
                when x"f1" & "0011" => d <= "00000000"; -- ........
                when x"f1" & "0100" => d <= "00011000"; -- ...##...
                when x"f1" & "0101" => d <= "00011000"; -- ...##...
                when x"f1" & "0110" => d <= "01111110"; -- .######.
                when x"f1" & "0111" => d <= "00011000"; -- ...##...
                when x"f1" & "1000" => d <= "00011000"; -- ...##...
                when x"f1" & "1001" => d <= "00000000"; -- ........
                when x"f1" & "1010" => d <= "00000000"; -- ........
                when x"f1" & "1011" => d <= "11111111"; -- ########
                when x"f1" & "1100" => d <= "00000000"; -- ........
                when x"f1" & "1101" => d <= "00000000"; -- ........
                when x"f1" & "1110" => d <= "00000000"; -- ........
                when x"f1" & "1111" => d <= "00000000"; -- ........

                when x"f2" & "0000" => d <= "00000000"; -- ........
                when x"f2" & "0001" => d <= "00000000"; -- ........
                when x"f2" & "0010" => d <= "00000000"; -- ........
                when x"f2" & "0011" => d <= "00110000"; -- ..##....
                when x"f2" & "0100" => d <= "00011000"; -- ...##...
                when x"f2" & "0101" => d <= "00001100"; -- ....##..
                when x"f2" & "0110" => d <= "00000110"; -- .....##.
                when x"f2" & "0111" => d <= "00001100"; -- ....##..
                when x"f2" & "1000" => d <= "00011000"; -- ...##...
                when x"f2" & "1001" => d <= "00110000"; -- ..##....
                when x"f2" & "1010" => d <= "00000000"; -- ........
                when x"f2" & "1011" => d <= "01111110"; -- .######.
                when x"f2" & "1100" => d <= "00000000"; -- ........
                when x"f2" & "1101" => d <= "00000000"; -- ........
                when x"f2" & "1110" => d <= "00000000"; -- ........
                when x"f2" & "1111" => d <= "00000000"; -- ........

                when x"f3" & "0000" => d <= "00000000"; -- ........
                when x"f3" & "0001" => d <= "00000000"; -- ........
                when x"f3" & "0010" => d <= "00000000"; -- ........
                when x"f3" & "0011" => d <= "00001100"; -- ....##..
                when x"f3" & "0100" => d <= "00011000"; -- ...##...
                when x"f3" & "0101" => d <= "00110000"; -- ..##....
                when x"f3" & "0110" => d <= "01100000"; -- .##.....
                when x"f3" & "0111" => d <= "00110000"; -- ..##....
                when x"f3" & "1000" => d <= "00011000"; -- ...##...
                when x"f3" & "1001" => d <= "00001100"; -- ....##..
                when x"f3" & "1010" => d <= "00000000"; -- ........
                when x"f3" & "1011" => d <= "01111110"; -- .######.
                when x"f3" & "1100" => d <= "00000000"; -- ........
                when x"f3" & "1101" => d <= "00000000"; -- ........
                when x"f3" & "1110" => d <= "00000000"; -- ........
                when x"f3" & "1111" => d <= "00000000"; -- ........

                when x"f4" & "0000" => d <= "00000000"; -- ........
                when x"f4" & "0001" => d <= "00000000"; -- ........
                when x"f4" & "0010" => d <= "00001110"; -- ....###.
                when x"f4" & "0011" => d <= "00011011"; -- ...##.##
                when x"f4" & "0100" => d <= "00011011"; -- ...##.##
                when x"f4" & "0101" => d <= "00011000"; -- ...##...
                when x"f4" & "0110" => d <= "00011000"; -- ...##...
                when x"f4" & "0111" => d <= "00011000"; -- ...##...
                when x"f4" & "1000" => d <= "00011000"; -- ...##...
                when x"f4" & "1001" => d <= "00011000"; -- ...##...
                when x"f4" & "1010" => d <= "00011000"; -- ...##...
                when x"f4" & "1011" => d <= "00011000"; -- ...##...
                when x"f4" & "1100" => d <= "00011000"; -- ...##...
                when x"f4" & "1101" => d <= "00011000"; -- ...##...
                when x"f4" & "1110" => d <= "00011000"; -- ...##...
                when x"f4" & "1111" => d <= "00011000"; -- ...##...

                when x"f5" & "0000" => d <= "00011000"; -- ...##...
                when x"f5" & "0001" => d <= "00011000"; -- ...##...
                when x"f5" & "0010" => d <= "00011000"; -- ...##...
                when x"f5" & "0011" => d <= "00011000"; -- ...##...
                when x"f5" & "0100" => d <= "00011000"; -- ...##...
                when x"f5" & "0101" => d <= "00011000"; -- ...##...
                when x"f5" & "0110" => d <= "00011000"; -- ...##...
                when x"f5" & "0111" => d <= "00011000"; -- ...##...
                when x"f5" & "1000" => d <= "11011000"; -- ##.##...
                when x"f5" & "1001" => d <= "11011000"; -- ##.##...
                when x"f5" & "1010" => d <= "11011000"; -- ##.##...
                when x"f5" & "1011" => d <= "01110000"; -- .###....
                when x"f5" & "1100" => d <= "00000000"; -- ........
                when x"f5" & "1101" => d <= "00000000"; -- ........
                when x"f5" & "1110" => d <= "00000000"; -- ........
                when x"f5" & "1111" => d <= "00000000"; -- ........

                when x"f6" & "0000" => d <= "00000000"; -- ........
                when x"f6" & "0001" => d <= "00000000"; -- ........
                when x"f6" & "0010" => d <= "00000000"; -- ........
                when x"f6" & "0011" => d <= "00000000"; -- ........
                when x"f6" & "0100" => d <= "00011000"; -- ...##...
                when x"f6" & "0101" => d <= "00011000"; -- ...##...
                when x"f6" & "0110" => d <= "00000000"; -- ........
                when x"f6" & "0111" => d <= "01111110"; -- .######.
                when x"f6" & "1000" => d <= "00000000"; -- ........
                when x"f6" & "1001" => d <= "00011000"; -- ...##...
                when x"f6" & "1010" => d <= "00011000"; -- ...##...
                when x"f6" & "1011" => d <= "00000000"; -- ........
                when x"f6" & "1100" => d <= "00000000"; -- ........
                when x"f6" & "1101" => d <= "00000000"; -- ........
                when x"f6" & "1110" => d <= "00000000"; -- ........
                when x"f6" & "1111" => d <= "00000000"; -- ........

                when x"f7" & "0000" => d <= "00000000"; -- ........
                when x"f7" & "0001" => d <= "00000000"; -- ........
                when x"f7" & "0010" => d <= "00000000"; -- ........
                when x"f7" & "0011" => d <= "00000000"; -- ........
                when x"f7" & "0100" => d <= "00000000"; -- ........
                when x"f7" & "0101" => d <= "01110110"; -- .###.##.
                when x"f7" & "0110" => d <= "11011100"; -- ##.###..
                when x"f7" & "0111" => d <= "00000000"; -- ........
                when x"f7" & "1000" => d <= "01110110"; -- .###.##.
                when x"f7" & "1001" => d <= "11011100"; -- ##.###..
                when x"f7" & "1010" => d <= "00000000"; -- ........
                when x"f7" & "1011" => d <= "00000000"; -- ........
                when x"f7" & "1100" => d <= "00000000"; -- ........
                when x"f7" & "1101" => d <= "00000000"; -- ........
                when x"f7" & "1110" => d <= "00000000"; -- ........
                when x"f7" & "1111" => d <= "00000000"; -- ........

                when x"f8" & "0000" => d <= "00000000"; -- ........
                when x"f8" & "0001" => d <= "00111000"; -- ..###...
                when x"f8" & "0010" => d <= "01101100"; -- .##.##..
                when x"f8" & "0011" => d <= "01101100"; -- .##.##..
                when x"f8" & "0100" => d <= "00111000"; -- ..###...
                when x"f8" & "0101" => d <= "00000000"; -- ........
                when x"f8" & "0110" => d <= "00000000"; -- ........
                when x"f8" & "0111" => d <= "00000000"; -- ........
                when x"f8" & "1000" => d <= "00000000"; -- ........
                when x"f8" & "1001" => d <= "00000000"; -- ........
                when x"f8" & "1010" => d <= "00000000"; -- ........
                when x"f8" & "1011" => d <= "00000000"; -- ........
                when x"f8" & "1100" => d <= "00000000"; -- ........
                when x"f8" & "1101" => d <= "00000000"; -- ........
                when x"f8" & "1110" => d <= "00000000"; -- ........
                when x"f8" & "1111" => d <= "00000000"; -- ........

                when x"f9" & "0000" => d <= "00000000"; -- ........
                when x"f9" & "0001" => d <= "00000000"; -- ........
                when x"f9" & "0010" => d <= "00000000"; -- ........
                when x"f9" & "0011" => d <= "00000000"; -- ........
                when x"f9" & "0100" => d <= "00000000"; -- ........
                when x"f9" & "0101" => d <= "00000000"; -- ........
                when x"f9" & "0110" => d <= "00000000"; -- ........
                when x"f9" & "0111" => d <= "00011000"; -- ...##...
                when x"f9" & "1000" => d <= "00011000"; -- ...##...
                when x"f9" & "1001" => d <= "00000000"; -- ........
                when x"f9" & "1010" => d <= "00000000"; -- ........
                when x"f9" & "1011" => d <= "00000000"; -- ........
                when x"f9" & "1100" => d <= "00000000"; -- ........
                when x"f9" & "1101" => d <= "00000000"; -- ........
                when x"f9" & "1110" => d <= "00000000"; -- ........
                when x"f9" & "1111" => d <= "00000000"; -- ........

                when x"fa" & "0000" => d <= "00000000"; -- ........
                when x"fa" & "0001" => d <= "00000000"; -- ........
                when x"fa" & "0010" => d <= "00000000"; -- ........
                when x"fa" & "0011" => d <= "00000000"; -- ........
                when x"fa" & "0100" => d <= "00000000"; -- ........
                when x"fa" & "0101" => d <= "00000000"; -- ........
                when x"fa" & "0110" => d <= "00000000"; -- ........
                when x"fa" & "0111" => d <= "00000000"; -- ........
                when x"fa" & "1000" => d <= "00011000"; -- ...##...
                when x"fa" & "1001" => d <= "00000000"; -- ........
                when x"fa" & "1010" => d <= "00000000"; -- ........
                when x"fa" & "1011" => d <= "00000000"; -- ........
                when x"fa" & "1100" => d <= "00000000"; -- ........
                when x"fa" & "1101" => d <= "00000000"; -- ........
                when x"fa" & "1110" => d <= "00000000"; -- ........
                when x"fa" & "1111" => d <= "00000000"; -- ........

                when x"fb" & "0000" => d <= "00000000"; -- ........
                when x"fb" & "0001" => d <= "00001111"; -- ....####
                when x"fb" & "0010" => d <= "00001100"; -- ....##..
                when x"fb" & "0011" => d <= "00001100"; -- ....##..
                when x"fb" & "0100" => d <= "00001100"; -- ....##..
                when x"fb" & "0101" => d <= "00001100"; -- ....##..
                when x"fb" & "0110" => d <= "00001100"; -- ....##..
                when x"fb" & "0111" => d <= "11101100"; -- ###.##..
                when x"fb" & "1000" => d <= "01101100"; -- .##.##..
                when x"fb" & "1001" => d <= "01101100"; -- .##.##..
                when x"fb" & "1010" => d <= "00111100"; -- ..####..
                when x"fb" & "1011" => d <= "00011100"; -- ...###..
                when x"fb" & "1100" => d <= "00000000"; -- ........
                when x"fb" & "1101" => d <= "00000000"; -- ........
                when x"fb" & "1110" => d <= "00000000"; -- ........
                when x"fb" & "1111" => d <= "00000000"; -- ........

                when x"fc" & "0000" => d <= "00000000"; -- ........
                when x"fc" & "0001" => d <= "11011000"; -- ##.##...
                when x"fc" & "0010" => d <= "01101100"; -- .##.##..
                when x"fc" & "0011" => d <= "01101100"; -- .##.##..
                when x"fc" & "0100" => d <= "01101100"; -- .##.##..
                when x"fc" & "0101" => d <= "01101100"; -- .##.##..
                when x"fc" & "0110" => d <= "01101100"; -- .##.##..
                when x"fc" & "0111" => d <= "00000000"; -- ........
                when x"fc" & "1000" => d <= "00000000"; -- ........
                when x"fc" & "1001" => d <= "00000000"; -- ........
                when x"fc" & "1010" => d <= "00000000"; -- ........
                when x"fc" & "1011" => d <= "00000000"; -- ........
                when x"fc" & "1100" => d <= "00000000"; -- ........
                when x"fc" & "1101" => d <= "00000000"; -- ........
                when x"fc" & "1110" => d <= "00000000"; -- ........
                when x"fc" & "1111" => d <= "00000000"; -- ........

                when x"fd" & "0000" => d <= "00000000"; -- ........
                when x"fd" & "0001" => d <= "01110000"; -- .###....
                when x"fd" & "0010" => d <= "11011000"; -- ##.##...
                when x"fd" & "0011" => d <= "00110000"; -- ..##....
                when x"fd" & "0100" => d <= "01100000"; -- .##.....
                when x"fd" & "0101" => d <= "11001000"; -- ##..#...
                when x"fd" & "0110" => d <= "11111000"; -- #####...
                when x"fd" & "0111" => d <= "00000000"; -- ........
                when x"fd" & "1000" => d <= "00000000"; -- ........
                when x"fd" & "1001" => d <= "00000000"; -- ........
                when x"fd" & "1010" => d <= "00000000"; -- ........
                when x"fd" & "1011" => d <= "00000000"; -- ........
                when x"fd" & "1100" => d <= "00000000"; -- ........
                when x"fd" & "1101" => d <= "00000000"; -- ........
                when x"fd" & "1110" => d <= "00000000"; -- ........
                when x"fd" & "1111" => d <= "00000000"; -- ........

                when x"fe" & "0000" => d <= "00000000"; -- ........
                when x"fe" & "0001" => d <= "00000000"; -- ........
                when x"fe" & "0010" => d <= "00000000"; -- ........
                when x"fe" & "0011" => d <= "00000000"; -- ........
                when x"fe" & "0100" => d <= "01111100"; -- .#####..
                when x"fe" & "0101" => d <= "01111100"; -- .#####..
                when x"fe" & "0110" => d <= "01111100"; -- .#####..
                when x"fe" & "0111" => d <= "01111100"; -- .#####..
                when x"fe" & "1000" => d <= "01111100"; -- .#####..
                when x"fe" & "1001" => d <= "01111100"; -- .#####..
                when x"fe" & "1010" => d <= "01111100"; -- .#####..
                when x"fe" & "1011" => d <= "00000000"; -- ........
                when x"fe" & "1100" => d <= "00000000"; -- ........
                when x"fe" & "1101" => d <= "00000000"; -- ........
                when x"fe" & "1110" => d <= "00000000"; -- ........
                when x"fe" & "1111" => d <= "00000000"; -- ........

                when x"ff" & "0000" => d <= "00000000"; -- ........
                when x"ff" & "0001" => d <= "00000000"; -- ........
                when x"ff" & "0010" => d <= "00000000"; -- ........
                when x"ff" & "0011" => d <= "00000000"; -- ........
                when x"ff" & "0100" => d <= "00000000"; -- ........
                when x"ff" & "0101" => d <= "00000000"; -- ........
                when x"ff" & "0110" => d <= "00000000"; -- ........
                when x"ff" & "0111" => d <= "00000000"; -- ........
                when x"ff" & "1000" => d <= "00000000"; -- ........
                when x"ff" & "1001" => d <= "00000000"; -- ........
                when x"ff" & "1010" => d <= "00000000"; -- ........
                when x"ff" & "1011" => d <= "00000000"; -- ........
                when x"ff" & "1100" => d <= "00000000"; -- ........
                when x"ff" & "1101" => d <= "00000000"; -- ........
                when x"ff" & "1110" => d <= "00000000"; -- ........
                when x"ff" & "1111" => d <= "00000000"; -- ........

                when others => d <= (others => '0');

            end case;
        end if;
    end process;

end architecture behavioural;
