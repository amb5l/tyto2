-- secure IP is supported by simulator, no substitution needed

configuration cfg_tb_hdmi_tpg of tb_hdmi_tpg is
  for sim
  end for;
end configuration cfg_tb_hdmi_tpg;
